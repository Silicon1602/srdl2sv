/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://github.com/Silicon1602/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : November 02 2021 23:27:37
 *  - Path     : /home/dpotter/srdl2sv/examples/enums
 *  - RDL file : ['enums.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : NONE
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Unpacked I/Os    : True
 *  - Register Bus Type: amba3ahblite
 *  - Address width    : 32
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': False, 'RegFile': False, 'Memory': False, 'Register': False, 'Field': False}
 *
 * ===LICENSE OF ENUMS.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module enums
    import enums_pkg::*;
    import enums__regfile_1_pkg::*;
(
    // Resets
     
    
    // Inputs
    input                                    clk                    ,
    input                                    HRESETn                ,
    input  [31:0]                            HADDR                  ,
    input                                    HWRITE                 ,
    input  [2:0]                             HSIZE                  ,
    input  [3:0]                             HPROT                  ,
    input  [1:0]                             HTRANS                 ,
    input  [32-1:0]                          HWDATA                 ,
    input                                    HSEL                   ,
    input  enums_pkg::third_enum             regfile_1__reg_c__f1_in,
    input  [1:0]                             regfile_1__reg_c__f2_in,
    input  enums__regfile_1_pkg::fourth_enum regfile_1__reg_d__f1_in,
    input  [1:0]                             regfile_1__reg_d__f2_in,
    input  enums_pkg::first_enum             reg_a__f1_in           ,
    input  [1:0]                             reg_a__f2_in           ,
    input  enums_pkg::second_enum            reg_b__f1_in           ,
    input  [1:0]                             reg_b__f2_in           ,
    
    // Outputs
    output                                   HREADYOUT             ,
    output                                   HRESP                 ,
    output [32-1:0]                          HRDATA                ,
    output enums_pkg::third_enum             regfile_1__reg_c__f1_r,
    output [1:0]                             regfile_1__reg_c__f2_r,
    output enums__regfile_1_pkg::fourth_enum regfile_1__reg_d__f1_r,
    output [1:0]                             regfile_1__reg_d__f2_r,
    output enums_pkg::first_enum             reg_a__f1_r           ,
    output [1:0]                             reg_a__f2_r           ,
    output enums_pkg::second_enum            reg_b__f1_r           ,
    output [1:0]                             reg_b__f2_r           
);


// Internal signals
srdl2sv_widget_if #(.ADDR_W (32), .DATA_W(32)) widget_if;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - widget_if -> SystemVerilog interface to between widgets
 *                   and the internal srdl2sv registers.
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA,

     // Interface to internal logic
     .widget_if);
/*******************************************************************
 *******************************************************************
 * REGFILE               : regfile_1
 * DIMENSION             : 0
 * DEPTHS (per dimension): []
 *******************************************************************
 *******************************************************************/


/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_c
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic                 regfile_1__reg_c_active     ;
logic                 regfile_1__reg_c_sw_wr      ;
logic [31:0]          regfile_1__reg_c_data_mux_in;
logic                 regfile_1__reg_c_rdy_mux_in ;
logic                 regfile_1__reg_c_err_mux_in ;
enums_pkg::third_enum regfile_1__reg_c__f1_q      ;
logic [1:0]           regfile_1__reg_c__f2_q      ;


// Register-activation for 'regfile_1__reg_c' 
assign regfile_1__reg_c_active = widget_if.addr == 8;
assign regfile_1__reg_c_sw_wr = regfile_1__reg_c_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (regfile_1__reg_c[1:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'encode']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_c_sw_wr)
    begin
        if (widget_if.byte_en[0])
            regfile_1__reg_c__f1_q[1:0] <= widget_if.w_data[1:0];
    end
    else
        // we or wel property not set
        regfile_1__reg_c__f1_q <= regfile_1__reg_c__f1_in;
end // of regfile_1__reg_c__f1's always_ff

// Connect register to hardware output port
assign regfile_1__reg_c__f1_r = regfile_1__reg_c__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (regfile_1__reg_c[9:8])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_c_sw_wr)
    begin
        if (widget_if.byte_en[1])
            regfile_1__reg_c__f2_q[1:0] <= widget_if.w_data[9:8];
    end
    else
        // we or wel property not set
        regfile_1__reg_c__f2_q <= regfile_1__reg_c__f2_in;
end // of regfile_1__reg_c__f2's always_ff

// Connect register to hardware output port
assign regfile_1__reg_c__f2_r = regfile_1__reg_c__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign regfile_1__reg_c_data_mux_in = {{22{1'b0}}, regfile_1__reg_c__f2_q, {6{1'b0}}, regfile_1__reg_c__f1_q};

// Internal registers are ready immediately
assign regfile_1__reg_c_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign regfile_1__reg_c_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_d
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic                             regfile_1__reg_d_active     ;
logic                             regfile_1__reg_d_sw_wr      ;
logic [31:0]                      regfile_1__reg_d_data_mux_in;
logic                             regfile_1__reg_d_rdy_mux_in ;
logic                             regfile_1__reg_d_err_mux_in ;
enums__regfile_1_pkg::fourth_enum regfile_1__reg_d__f1_q      ;
logic [1:0]                       regfile_1__reg_d__f2_q      ;


// Register-activation for 'regfile_1__reg_d' 
assign regfile_1__reg_d_active = widget_if.addr == 12;
assign regfile_1__reg_d_sw_wr = regfile_1__reg_d_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (regfile_1__reg_d[1:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'encode']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_d_sw_wr)
    begin
        if (widget_if.byte_en[0])
            regfile_1__reg_d__f1_q[1:0] <= widget_if.w_data[1:0];
    end
    else
        // we or wel property not set
        regfile_1__reg_d__f1_q <= regfile_1__reg_d__f1_in;
end // of regfile_1__reg_d__f1's always_ff

// Connect register to hardware output port
assign regfile_1__reg_d__f1_r = regfile_1__reg_d__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (regfile_1__reg_d[9:8])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_d_sw_wr)
    begin
        if (widget_if.byte_en[1])
            regfile_1__reg_d__f2_q[1:0] <= widget_if.w_data[9:8];
    end
    else
        // we or wel property not set
        regfile_1__reg_d__f2_q <= regfile_1__reg_d__f2_in;
end // of regfile_1__reg_d__f2's always_ff

// Connect register to hardware output port
assign regfile_1__reg_d__f2_r = regfile_1__reg_d__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign regfile_1__reg_d_data_mux_in = {{22{1'b0}}, regfile_1__reg_d__f2_q, {6{1'b0}}, regfile_1__reg_d__f1_q};

// Internal registers are ready immediately
assign regfile_1__reg_d_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign regfile_1__reg_d_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_a
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic                 reg_a_active     ;
logic                 reg_a_sw_wr      ;
logic [31:0]          reg_a_data_mux_in;
logic                 reg_a_rdy_mux_in ;
logic                 reg_a_err_mux_in ;
enums_pkg::first_enum reg_a__f1_q      ;
logic [1:0]           reg_a__f2_q      ;


// Register-activation for 'reg_a' 
assign reg_a_active = widget_if.addr == 0;
assign reg_a_sw_wr = reg_a_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (reg_a[1:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'encode']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_a_sw_wr)
    begin
        if (widget_if.byte_en[0])
            reg_a__f1_q[1:0] <= widget_if.w_data[1:0];
    end
    else
        // we or wel property not set
        reg_a__f1_q <= reg_a__f1_in;
end // of reg_a__f1's always_ff

// Connect register to hardware output port
assign reg_a__f1_r = reg_a__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (reg_a[9:8])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_a_sw_wr)
    begin
        if (widget_if.byte_en[1])
            reg_a__f2_q[1:0] <= widget_if.w_data[9:8];
    end
    else
        // we or wel property not set
        reg_a__f2_q <= reg_a__f2_in;
end // of reg_a__f2's always_ff

// Connect register to hardware output port
assign reg_a__f2_r = reg_a__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg_a_data_mux_in = {{22{1'b0}}, reg_a__f2_q, {6{1'b0}}, reg_a__f1_q};

// Internal registers are ready immediately
assign reg_a_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg_a_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_b
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic                  reg_b_active     ;
logic                  reg_b_sw_wr      ;
logic [31:0]           reg_b_data_mux_in;
logic                  reg_b_rdy_mux_in ;
logic                  reg_b_err_mux_in ;
enums_pkg::second_enum reg_b__f1_q      ;
logic [1:0]            reg_b__f2_q      ;


// Register-activation for 'reg_b' 
assign reg_b_active = widget_if.addr == 4;
assign reg_b_sw_wr = reg_b_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (reg_b[1:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'encode']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_b_sw_wr)
    begin
        if (widget_if.byte_en[0])
            reg_b__f1_q[1:0] <= widget_if.w_data[1:0];
    end
    else
        // we or wel property not set
        reg_b__f1_q <= reg_b__f1_in;
end // of reg_b__f1's always_ff

// Connect register to hardware output port
assign reg_b__f1_r = reg_b__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (reg_b[9:8])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_b_sw_wr)
    begin
        if (widget_if.byte_en[1])
            reg_b__f2_q[1:0] <= widget_if.w_data[9:8];
    end
    else
        // we or wel property not set
        reg_b__f2_q <= reg_b__f2_in;
end // of reg_b__f2's always_ff

// Connect register to hardware output port
assign reg_b__f2_r = reg_b__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg_b_data_mux_in = {{22{1'b0}}, reg_b__f2_q, {6{1'b0}}, reg_b__f1_q};

// Internal registers are ready immediately
assign reg_b_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg_b_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0])));

// Read multiplexer
always_comb
begin
    unique case (1'b1)
        regfile_1__reg_c_active:
        begin
            widget_if.r_data = regfile_1__reg_c_data_mux_in;
            widget_if.err    = regfile_1__reg_c_err_mux_in;
            widget_if.rdy    = regfile_1__reg_c_rdy_mux_in;
        end
        regfile_1__reg_d_active:
        begin
            widget_if.r_data = regfile_1__reg_d_data_mux_in;
            widget_if.err    = regfile_1__reg_d_err_mux_in;
            widget_if.rdy    = regfile_1__reg_d_rdy_mux_in;
        end
        reg_a_active:
        begin
            widget_if.r_data = reg_a_data_mux_in;
            widget_if.err    = reg_a_err_mux_in;
            widget_if.rdy    = reg_a_rdy_mux_in;
        end
        reg_b_active:
        begin
            widget_if.r_data = reg_b_data_mux_in;
            widget_if.err    = reg_b_err_mux_in;
            widget_if.rdy    = reg_b_rdy_mux_in;
        end
        default:
        begin
            // If the address is not found, return an error
            widget_if.r_data = 0;
            widget_if.err    = 1;
            widget_if.rdy    = widget_if.r_vld || widget_if.w_vld;
        end
    endcase
end
endmodule
