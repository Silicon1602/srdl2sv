/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://github.com/Silicon1602/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : November 07 2021 11:16:51
 *  - Path     : /home/dpotter/srdl2sv/examples/aliases
 *  - RDL file : ['aliases.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : NONE
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Address Errors   : True
 *  - Unpacked I/Os    : True
 *  - Register Bus Type: amba3ahblite
 *  - Address width    : 32
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': True, 'RegFile': True, 'Memory': True, 'Register': True, 'Field': True}
 *
 * ===LICENSE OF ALIASES.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module aliases
    
(
    // Resets
     
    
    // Inputs
    input               clk                                    ,
    input               HRESETn                                ,
    input  [31:0]       HADDR                                  ,
    input               HWRITE                                 ,
    input  [2:0]        HSIZE                                  ,
    input  [3:0]        HPROT                                  ,
    input  [1:0]        HTRANS                                 ,
    input  [32-1:0]     HWDATA                                 ,
    input               HSEL                                   ,
    input               example_rf__ext_main_reg__f1_ext_r_err [4],
    input               example_rf__ext_main_reg__f1_ext_r_ack [4],
    input               example_rf__ext_main_reg__f2_ext_r_err [4],
    input               example_rf__ext_main_reg__f2_ext_r_ack [4],
    input               example_rf__ext_main_reg__f1_ext_w_err [4],
    input               example_rf__ext_main_reg__f1_ext_w_ack [4],
    input               example_rf__ext_main_reg__f2_ext_w_err [4],
    input               example_rf__ext_main_reg__f2_ext_w_ack [4],
    input  [15:0]       example_rf__ext_main_reg__f1_ext_r_data[4],
    input  [15:0]       example_rf__ext_main_reg__f2_ext_r_data[4],
    input  [0:0]        event1__some_event_in                  ,
    input               four_field_reg__f1_hw_wr               ,
    input  [7:0]        four_field_reg__f1_in                  ,
    input               four_field_reg__f2_hw_wr               ,
    input  [7:0]        four_field_reg__f2_in                  ,
    input               four_field_reg__f3_hw_wr               ,
    input  [7:0]        four_field_reg__f3_in                  ,
    input               four_field_reg__f4_hw_wr               ,
    input  [7:0]        four_field_reg__f4_in                  ,
    
    // Outputs
    output              HREADYOUT                               ,
    output              HRESP                                   ,
    output [32-1:0]     HRDATA                                  ,
    output              example_rf__ext_main_reg__f1_ext_w_req  [4],
    output [15:0]       example_rf__ext_main_reg__f1_ext_w_data [4],
    output [15:0]       example_rf__ext_main_reg__f1_ext_w_mask [4],
    output              example_rf__ext_main_reg__f1_ext_r_req  [4],
    output              example_rf__ext_alias_reg__field_1_ext_w_req[4],
    output [15:0]       example_rf__ext_alias_reg__field_1_ext_w_data[4],
    output [15:0]       example_rf__ext_alias_reg__field_1_ext_w_mask[4],
    output              example_rf__ext_alias_reg__field_1_ext_r_req[4],
    output              example_rf__ext_main_reg__f2_ext_w_req  [4],
    output [15:0]       example_rf__ext_main_reg__f2_ext_w_data [4],
    output [15:0]       example_rf__ext_main_reg__f2_ext_w_mask [4],
    output              example_rf__ext_main_reg__f2_ext_r_req  [4],
    output              event1_intr                             ,
    output [7:0]        four_field_reg__f1_r                    ,
    output [7:0]        four_field_reg__f2_r                    ,
    output [7:0]        four_field_reg__f3_r                    ,
    output reg          four_field_reg__f3_swmod                ,
    output [7:0]        four_field_reg__f4_r                    
);


// Internal signals
srdl2sv_widget_if #(.ADDR_W (32), .DATA_W(32)) widget_if;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - widget_if -> SystemVerilog interface to between widgets
 *                   and the internal srdl2sv registers.
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA,

     // Interface to internal logic
     .widget_if);

genvar gv_a;

/*******************************************************************
 *******************************************************************
 * REGFILE               : example_rf
 * DIMENSION             : 1
 * DEPTHS (per dimension): [4]
 *******************************************************************
 *******************************************************************/

/**REGFILE DESCRIPTION**********************************************
Instantiate regfile to show that they also work in regfiles.
/*******************************************************************/

// Variables of register 'ext_main_reg'
logic        example_rf__ext_main_reg_active      [4];
logic        example_rf__ext_main_reg_sw_rd       [4];
logic        example_rf__ext_main_reg_sw_wr       [4];
logic        example_rf__ext_alias_reg_active     [4];
logic        example_rf__ext_alias_reg_sw_rd      [4];
logic        example_rf__ext_alias_reg_sw_wr      [4];
logic [31:0] example_rf__ext_main_reg_data_mux_in [4];
logic        example_rf__ext_main_reg_rdy_mux_in  [4];
logic        example_rf__ext_main_reg_err_mux_in  [4];
logic [31:0] example_rf__ext_alias_reg_data_mux_in[4];
logic        example_rf__ext_alias_reg_rdy_mux_in [4];
logic        example_rf__ext_alias_reg_err_mux_in [4];
logic [15:0] example_rf__ext_main_reg__f1_q       [4];
logic [15:0] example_rf__ext_alias_reg__field_1_q [4];
logic [15:0] example_rf__ext_main_reg__f2_q       [4];

generate
for (gv_a = 0; gv_a < 4; gv_a++)
begin
    
    /*******************************************************************
    /*******************************************************************
    /* REGISTER              : ext_main_reg
    /* DIMENSION             : 0
    /* DEPTHS (per dimension): []
    /*******************************************************************
    /*******************************************************************/
    
    /**REGISTER DESCRIPTION*********************************************
    If aliases registers are declared to be external,
    the external hardware will get a seperate interface
    for those registers.
    /*******************************************************************/
    
    // Register-activation for 'example_rf__ext_main_reg' 
    assign example_rf__ext_main_reg_active[gv_a] = widget_if.addr == 16+(gv_a*8);
    assign example_rf__ext_main_reg_sw_rd[gv_a] = example_rf__ext_main_reg_active[gv_a] && widget_if.r_vld;
    assign example_rf__ext_main_reg_sw_wr[gv_a] = example_rf__ext_main_reg_active[gv_a] && widget_if.w_vld;
    
    // Register-activation for 'example_rf__ext_alias_reg' (alias)
    assign example_rf__ext_alias_reg_active[gv_a] = widget_if.addr == 20+(gv_a*8);
    assign example_rf__ext_alias_reg_sw_rd[gv_a] = example_rf__ext_alias_reg_active[gv_a] && widget_if.r_vld;
    assign example_rf__ext_alias_reg_sw_wr[gv_a] = example_rf__ext_alias_reg_active[gv_a] && widget_if.w_vld;
    
    //-----------------FIELD SUMMARY-----------------
    // name         : f1 (example_rf__ext_main_reg[15:0])
    // access       : hw = rw  
    //                sw = rw (precedence)
    // reset        : - / -
    // flags        : ['sw', 'wel']
    // external     : True
    // storage type : StorageType.FLOPS
    //-----------------------------------------------
    
    
    /***********************************
     * Handle external write interface *
     ***********************************
     * The 'example_rf__ext_main_reg__f1_ext_w_req' output will be asserted once a write
     * is requested by the bus and will stay high until 'example_rf__ext_main_reg__f1_ext_w_ack' 
     * gets set. During a write, hardware shall not touch any bits that
     * are not defined in 'example_rf__ext_main_reg__f1_ext_w_mask'.
     *
     * 'example_rf__ext_main_reg__f1_ext_w_ack' shall be held 1'b1 until all fields in the register
     * acknowledged the read. In practice, this means until 'example_rf__ext_main_reg__f1_ext_w_req'
     * goes back to 1'b0.
     *
     * If 'example_rf__ext_main_reg__f1_ext_w_err' gets set, it must also be held during the
     * complete time 'example_rf__ext_main_reg__f1_ext_w_ack' is high.
     */
    // Write request
    assign example_rf__ext_main_reg__f1_ext_w_req[gv_a] = example_rf__ext_main_reg_sw_wr[gv_a];
    
    // Assign value from bus to output
    assign example_rf__ext_main_reg__f1_ext_w_data[gv_a] = widget_if.w_data[15:0];
    
    // Provide bit-wise mask. Only bits set to 1'b1 shall be written
    assign example_rf__ext_main_reg__f1_ext_w_mask[gv_a] = {{8{widget_if.byte_en[1]}},{8{widget_if.byte_en[0]}}};
    
    /**********************************
     * Handle external read interface *
     **********************************
     * The 'example_rf__ext_main_reg__f1_ext_r_req' output will be asserted once a read
     * is requested by the bus and will stay high until 'example_rf__ext_main_reg__f1_ext_r_ack' 
     * gets set. During a read, byte-enables will be ignored.
     *
     * 'example_rf__ext_main_reg__f1_ext_r_ack' shall be held 1'b1 until all fields in the register
     * acknowledged the read. In practice, this means until 'example_rf__ext_main_reg__f1_ext_r_req'
     * goes back to 1'b0.
     *
     * If 'example_rf__ext_main_reg__f1_ext_r_err' gets set, it must also be held during the
     * complete time 'example_rf__ext_main_reg__f1_ext_r_ack' is high.
     */
    // Actual data
    assign example_rf__ext_main_reg__f1_ext_r_req[gv_a] = example_rf__ext_main_reg_sw_rd[gv_a];
    
    // Assign return from outside hardware
    assign example_rf__ext_main_reg__f1_q[gv_a] = example_rf__ext_main_reg__f1_ext_r_data;
    
    /**********************************
     * Alias external write interface *
     **********************************
     * The hardware gets notified via a different wire that 
     * software accessed the register via an alias, but the return
     * shall be done via the main register's I/O. This is similar to
     * the implementation of an alias registers.
     */
    assign example_rf__ext_alias_reg__field_1_ext_w_req[gv_a] = example_rf__ext_alias_reg_sw_wr[gv_a];
    assign example_rf__ext_alias_reg__field_1_ext_w_data[gv_a] = widget_if.w_data[15:0];
    assign example_rf__ext_alias_reg__field_1_ext_w_mask[gv_a] = {{8{widget_if.byte_en[1]}},{8{widget_if.byte_en[0]}}};
    
    /*********************************
     * Alias external read interface *
     *********************************
     * The hardware gets notified via a different wire that 
     * software accessed the register via an alias, but the return
     * shall be done via the main register's I/O. This is similar to
     * the implementation of an alias registers.
     */
    assign example_rf__ext_alias_reg__field_1_ext_r_req[gv_a] = example_rf__ext_alias_reg_sw_rd[gv_a];
    
    //-----------------FIELD SUMMARY-----------------
    // name         : f2 (example_rf__ext_main_reg[31:16])
    // access       : hw = rw  
    //                sw = rw (precedence)
    // reset        : - / -
    // flags        : ['sw', 'wel']
    // external     : True
    // storage type : StorageType.FLOPS
    //-----------------------------------------------
    
    
    /***********************************
     * Handle external write interface *
     ***********************************
     * The 'example_rf__ext_main_reg__f2_ext_w_req' output will be asserted once a write
     * is requested by the bus and will stay high until 'example_rf__ext_main_reg__f2_ext_w_ack' 
     * gets set. During a write, hardware shall not touch any bits that
     * are not defined in 'example_rf__ext_main_reg__f2_ext_w_mask'.
     *
     * 'example_rf__ext_main_reg__f2_ext_w_ack' shall be held 1'b1 until all fields in the register
     * acknowledged the read. In practice, this means until 'example_rf__ext_main_reg__f2_ext_w_req'
     * goes back to 1'b0.
     *
     * If 'example_rf__ext_main_reg__f2_ext_w_err' gets set, it must also be held during the
     * complete time 'example_rf__ext_main_reg__f2_ext_w_ack' is high.
     */
    // Write request
    assign example_rf__ext_main_reg__f2_ext_w_req[gv_a] = example_rf__ext_main_reg_sw_wr[gv_a];
    
    // Assign value from bus to output
    assign example_rf__ext_main_reg__f2_ext_w_data[gv_a] = widget_if.w_data[31:16];
    
    // Provide bit-wise mask. Only bits set to 1'b1 shall be written
    assign example_rf__ext_main_reg__f2_ext_w_mask[gv_a] = {{8{widget_if.byte_en[3]}},{8{widget_if.byte_en[2]}}};
    
    /**********************************
     * Handle external read interface *
     **********************************
     * The 'example_rf__ext_main_reg__f2_ext_r_req' output will be asserted once a read
     * is requested by the bus and will stay high until 'example_rf__ext_main_reg__f2_ext_r_ack' 
     * gets set. During a read, byte-enables will be ignored.
     *
     * 'example_rf__ext_main_reg__f2_ext_r_ack' shall be held 1'b1 until all fields in the register
     * acknowledged the read. In practice, this means until 'example_rf__ext_main_reg__f2_ext_r_req'
     * goes back to 1'b0.
     *
     * If 'example_rf__ext_main_reg__f2_ext_r_err' gets set, it must also be held during the
     * complete time 'example_rf__ext_main_reg__f2_ext_r_ack' is high.
     */
    // Actual data
    assign example_rf__ext_main_reg__f2_ext_r_req[gv_a] = example_rf__ext_main_reg_sw_rd[gv_a];
    
    // Assign return from outside hardware
    assign example_rf__ext_main_reg__f2_q[gv_a] = example_rf__ext_main_reg__f2_ext_r_data;
    
    
    /********************************************** 
     * Assign all fields to signal to Mux         *
     **********************************************/
    // Assign all fields. Fields that are not readable are tied to 0.
    assign example_rf__ext_main_reg_data_mux_in[gv_a] = {example_rf__ext_main_reg__f2_q[gv_a], example_rf__ext_main_reg__f1_q[gv_a]};
    
    // Internal registers are ready immediately
    assign example_rf__ext_main_reg_rdy_mux_in[gv_a] = (example_rf__ext_main_reg__f1_ext_r_ack[gv_a] && example_rf__ext_main_reg__f2_ext_r_ack[gv_a] && widget_if.r_vld) || (example_rf__ext_main_reg__f1_ext_w_ack[gv_a] && example_rf__ext_main_reg__f2_ext_w_ack[gv_a] && widget_if.w_vld);
    
    // Return an error if *no* read and *no* write was succesful. If some bits
    // cannot be read/written but others are succesful, don't return and error
    // Hence, as long as one action can be succesful, no error will be returned.
    assign example_rf__ext_main_reg_err_mux_in[gv_a] = !((widget_if.r_vld && (|widget_if.byte_en[3:0])) || (widget_if.w_vld && (|widget_if.byte_en[3:0]))) || (example_rf__ext_main_reg__f1_ext_r_err[gv_a] && example_rf__ext_main_reg__f1_ext_r_ack[gv_a] && widget_if.r_vld) || (example_rf__ext_main_reg__f2_ext_r_err[gv_a] && example_rf__ext_main_reg__f2_ext_r_ack[gv_a] && widget_if.r_vld) || (example_rf__ext_main_reg__f1_ext_w_err[gv_a] && example_rf__ext_main_reg__f1_ext_w_ack[gv_a] && widget_if.w_vld) || (example_rf__ext_main_reg__f2_ext_w_err[gv_a] && example_rf__ext_main_reg__f2_ext_w_ack[gv_a] && widget_if.w_vld);
    
    /********************************************** 
     * Assign all fields to signal to Mux (alias) *
     **********************************************/
    // Assign all fields. Fields that are not readable are tied to 0.
    assign example_rf__ext_alias_reg_data_mux_in[gv_a] = {{16{1'b0}}, example_rf__ext_main_reg__f1_q[gv_a]};
    
    // Internal registers are ready immediately
    assign example_rf__ext_alias_reg_rdy_mux_in[gv_a] = (example_rf__ext_main_reg__f1_ext_r_ack[gv_a] && example_rf__ext_main_reg__f2_ext_r_ack[gv_a] && widget_if.r_vld) || (example_rf__ext_main_reg__f1_ext_w_ack[gv_a] && example_rf__ext_main_reg__f2_ext_w_ack[gv_a] && widget_if.w_vld);
    
    // Return an error if *no* read and *no* write was succesful. If some bits
    // cannot be read/written but others are succesful, don't return and error
    // Hence, as long as one action can be succesful, no error will be returned.
    assign example_rf__ext_alias_reg_err_mux_in[gv_a] = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0]))) || (example_rf__ext_main_reg__f1_ext_r_err[gv_a] && example_rf__ext_main_reg__f1_ext_r_ack[gv_a] && widget_if.r_vld) || (example_rf__ext_main_reg__f1_ext_w_err[gv_a] && example_rf__ext_main_reg__f1_ext_w_ack[gv_a] && widget_if.w_vld);
end // of for loop with iterator gv_a
endgenerate


/*******************************************************************
/*******************************************************************
/* REGISTER              : event1
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

/**REGISTER DESCRIPTION*********************************************
This register shows the alias example from Section 10.5.2 of the
SystemRDL2.0 spec (with some slight adaptations to make it compilable).
/*******************************************************************/
logic        event1_active                  ;
logic        event1_sw_wr                   ;
logic        event1_for_dv_active           ;
logic        event1_for_dv_sw_wr            ;
logic [31:0] event1_data_mux_in             ;
logic        event1_rdy_mux_in              ;
logic        event1_err_mux_in              ;
logic [31:0] event1_for_dv_data_mux_in      ;
logic        event1_for_dv_rdy_mux_in       ;
logic        event1_for_dv_err_mux_in       ;
logic [0:0]  event1__some_event_sticky_latch;
logic [0:0]  event1__some_event_q           ;


// Register-activation for 'event1' 
assign event1_active = widget_if.addr == 0;
assign event1_sw_wr = event1_active && widget_if.w_vld;

// Register-activation for 'event1_for_dv' (alias)
assign event1_for_dv_active = widget_if.addr == 4;
assign event1_for_dv_sw_wr = event1_for_dv_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : some_event (event1[0:0])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['intr', 'intr type', 'sw', 'woclr']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (event1_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
            event1__some_event_q[0:0] <= event1__some_event_q[0:0] & ~widget_if.w_data[0:0];
    end
    else
    if (event1_for_dv_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woset property
            event1__some_event_q[0:0] <= event1__some_event_q[0:0] | widget_if.w_data[0:0];
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (event1__some_event_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                event1__some_event_q[i] <= 1'b1;
            end
        end
    end
end // of event1__some_event's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign event1__some_event_sticky_latch = event1__some_event_in;


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign event1_intr = |(event1__some_event_q);


/********************************************** 
 * Assign all fields to signal to Mux         *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign event1_data_mux_in = {{31{1'b0}}, event1__some_event_q};

// Internal registers are ready immediately
assign event1_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign event1_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/********************************************** 
 * Assign all fields to signal to Mux (alias) *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign event1_for_dv_data_mux_in = {{31{1'b0}}, event1__some_event_q};

// Internal registers are ready immediately
assign event1_for_dv_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign event1_for_dv_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : four_field_reg
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

/**REGISTER DESCRIPTION*********************************************
This is a register with 4 fields.
/*******************************************************************/
logic        four_field_reg_active          ;
logic        four_field_reg_sw_wr           ;
logic        two_field_alias_active         ;
logic        two_field_alias_sw_wr          ;
logic        four_field_reg__any_alias_sw_wr;
logic [31:0] four_field_reg_data_mux_in     ;
logic        four_field_reg_rdy_mux_in      ;
logic        four_field_reg_err_mux_in      ;
logic [31:0] two_field_alias_data_mux_in    ;
logic        two_field_alias_rdy_mux_in     ;
logic        two_field_alias_err_mux_in     ;
logic [7:0]  four_field_reg__f1_q           ;
logic [7:0]  four_field_reg__f2_q           ;
logic [7:0]  four_field_reg__f3_q           ;
logic [7:0]  four_field_reg__f4_q           ;


// Register-activation for 'four_field_reg' 
assign four_field_reg_active = widget_if.addr == 8;
assign four_field_reg_sw_wr = four_field_reg_active && widget_if.w_vld;

// Register-activation for 'two_field_alias' (alias)
assign two_field_alias_active = widget_if.addr == 12;
assign two_field_alias_sw_wr = two_field_alias_active && widget_if.w_vld;

// Combined register activation. These will become active on
// access via any of the alias registers.
assign four_field_reg__any_alias_sw_wr = four_field_reg_sw_wr || two_field_alias_sw_wr;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (four_field_reg[7:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'wel']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (four_field_reg_sw_wr)
    begin
        if (widget_if.byte_en[0])
            four_field_reg__f1_q[7:0] <= widget_if.w_data[7:0];
    end
    else
    if (two_field_alias_sw_wr)
    begin
        if (widget_if.byte_en[0])
            four_field_reg__f1_q[7:0] <= widget_if.w_data[7:0];
    end
    else
    if (!four_field_reg__f1_hw_wr)
        four_field_reg__f1_q <= four_field_reg__f1_in;
end // of four_field_reg__f1's always_ff

// Connect register to hardware output port
assign four_field_reg__f1_r = four_field_reg__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (four_field_reg[15:8])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'wel']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (four_field_reg_sw_wr)
    begin
        if (widget_if.byte_en[1])
            four_field_reg__f2_q[7:0] <= widget_if.w_data[15:8];
    end
    else
    if (!four_field_reg__f2_hw_wr)
        four_field_reg__f2_q <= four_field_reg__f2_in;
end // of four_field_reg__f2's always_ff

// Connect register to hardware output port
assign four_field_reg__f2_r = four_field_reg__f2_q;



//-----------------FIELD SUMMARY-----------------
// name         : f3 (four_field_reg[23:16])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'wel', 'swmod']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (four_field_reg_sw_wr)
    begin
        if (widget_if.byte_en[2])
            four_field_reg__f3_q[7:0] <= widget_if.w_data[23:16];
    end
    else
    if (!four_field_reg__f3_hw_wr)
        four_field_reg__f3_q <= four_field_reg__f3_in;
end // of four_field_reg__f3's always_ff

// Connect register to hardware output port
assign four_field_reg__f3_r = four_field_reg__f3_q;

// Combinational block to generate swmod-output signals
always_comb
begin
    four_field_reg__f3_swmod  = 0;
    four_field_reg__f3_swmod |= four_field_reg__any_alias_sw_wr && |widget_if.byte_en[2:2];
end


//-----------------FIELD SUMMARY-----------------
// name         : f4 (four_field_reg[31:24])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'wel', 'rclr']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (four_field_reg_sw_wr)
    begin
        if (widget_if.byte_en[3])
            four_field_reg__f4_q[7:0] <= widget_if.w_data[31:24];
    end
    else
    if (two_field_alias_sw_wr)
    begin
        if (widget_if.byte_en[3]) // woclr property
            four_field_reg__f4_q[7:0] <= four_field_reg__f4_q[7:0] & ~widget_if.w_data[31:24];
    end
    else
    if (!four_field_reg__f4_hw_wr)
        four_field_reg__f4_q <= four_field_reg__f4_in;
end // of four_field_reg__f4's always_ff

// Connect register to hardware output port
assign four_field_reg__f4_r = four_field_reg__f4_q;




/********************************************** 
 * Assign all fields to signal to Mux         *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign four_field_reg_data_mux_in = {four_field_reg__f4_q, four_field_reg__f3_q, four_field_reg__f2_q, four_field_reg__f1_q};

// Internal registers are ready immediately
assign four_field_reg_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign four_field_reg_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[3:0])) || (widget_if.w_vld && (|widget_if.byte_en[3:0])));

/********************************************** 
 * Assign all fields to signal to Mux (alias) *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign two_field_alias_data_mux_in = {four_field_reg__f4_q, {16{1'b0}}, four_field_reg__f1_q};

// Internal registers are ready immediately
assign two_field_alias_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign two_field_alias_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[3] || widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[3] || widget_if.byte_en[0])));

// Read multiplexer
always_comb
begin
    unique case (1'b1)
        example_rf__ext_main_reg_active[0]:
        begin
            widget_if.r_data = example_rf__ext_main_reg_data_mux_in[0];
            widget_if.err    = example_rf__ext_main_reg_err_mux_in[0];
            widget_if.rdy    = example_rf__ext_main_reg_rdy_mux_in[0];
        end
        example_rf__ext_main_reg_active[1]:
        begin
            widget_if.r_data = example_rf__ext_main_reg_data_mux_in[1];
            widget_if.err    = example_rf__ext_main_reg_err_mux_in[1];
            widget_if.rdy    = example_rf__ext_main_reg_rdy_mux_in[1];
        end
        example_rf__ext_main_reg_active[2]:
        begin
            widget_if.r_data = example_rf__ext_main_reg_data_mux_in[2];
            widget_if.err    = example_rf__ext_main_reg_err_mux_in[2];
            widget_if.rdy    = example_rf__ext_main_reg_rdy_mux_in[2];
        end
        example_rf__ext_main_reg_active[3]:
        begin
            widget_if.r_data = example_rf__ext_main_reg_data_mux_in[3];
            widget_if.err    = example_rf__ext_main_reg_err_mux_in[3];
            widget_if.rdy    = example_rf__ext_main_reg_rdy_mux_in[3];
        end
        example_rf__ext_alias_reg_active[0]:
        begin
            widget_if.r_data = example_rf__ext_alias_reg_data_mux_in[0];
            widget_if.err    = example_rf__ext_alias_reg_err_mux_in[0];
            widget_if.rdy    = example_rf__ext_alias_reg_rdy_mux_in[0];
        end
        example_rf__ext_alias_reg_active[1]:
        begin
            widget_if.r_data = example_rf__ext_alias_reg_data_mux_in[1];
            widget_if.err    = example_rf__ext_alias_reg_err_mux_in[1];
            widget_if.rdy    = example_rf__ext_alias_reg_rdy_mux_in[1];
        end
        example_rf__ext_alias_reg_active[2]:
        begin
            widget_if.r_data = example_rf__ext_alias_reg_data_mux_in[2];
            widget_if.err    = example_rf__ext_alias_reg_err_mux_in[2];
            widget_if.rdy    = example_rf__ext_alias_reg_rdy_mux_in[2];
        end
        example_rf__ext_alias_reg_active[3]:
        begin
            widget_if.r_data = example_rf__ext_alias_reg_data_mux_in[3];
            widget_if.err    = example_rf__ext_alias_reg_err_mux_in[3];
            widget_if.rdy    = example_rf__ext_alias_reg_rdy_mux_in[3];
        end
        event1_active:
        begin
            widget_if.r_data = event1_data_mux_in;
            widget_if.err    = event1_err_mux_in;
            widget_if.rdy    = event1_rdy_mux_in;
        end
        event1_for_dv_active:
        begin
            widget_if.r_data = event1_for_dv_data_mux_in;
            widget_if.err    = event1_for_dv_err_mux_in;
            widget_if.rdy    = event1_for_dv_rdy_mux_in;
        end
        four_field_reg_active:
        begin
            widget_if.r_data = four_field_reg_data_mux_in;
            widget_if.err    = four_field_reg_err_mux_in;
            widget_if.rdy    = four_field_reg_rdy_mux_in;
        end
        two_field_alias_active:
        begin
            widget_if.r_data = two_field_alias_data_mux_in;
            widget_if.err    = two_field_alias_err_mux_in;
            widget_if.rdy    = two_field_alias_rdy_mux_in;
        end
        default:
        begin
            // If the address is not found, return an error
            widget_if.r_data = 0;
            widget_if.err    = 1;
            widget_if.rdy    = widget_if.r_vld || widget_if.w_vld;
        end
    endcase
end
endmodule
