/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://github.com/Silicon1602/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : November 26 2021 16:33:16
 *  - Path     : /home/dpotter/srdl2sv/examples/parameters
 *  - RDL file : ['parameters.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : NONE
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Address Errors   : True
 *  - Unpacked I/Os    : True
 *  - Register Bus Type: amba3ahblite
 *  - Address width    : 32
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': False, 'RegFile': False, 'Memory': False, 'Register': False, 'Field': False}
 *
 * ===LICENSE OF PAREMETERS.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module paremeters
    
(
    // Reset signals declared for registers
    input  rst_async_n, 
    
    // Ports for 'General Clock'
    input               clk,
    
    // Ports for 'AHB Protocol'
    input               HRESETn  ,
    input  [31:0]       HADDR    ,
    input               HWRITE   ,
    input  [2:0]        HSIZE    ,
    input  [3:0]        HPROT    ,
    input  [1:0]        HTRANS   ,
    input  [32-1:0]     HWDATA   ,
    input               HSEL     ,
    output              HREADYOUT,
    output              HRESP    ,
    output [32-1:0]     HRDATA   ,
    
    // Ports for 'reg32'
    input  [31:0]       reg32__data_in,
    output [31:0]       reg32__data_r ,
    
    // Ports for 'reg32_arr'
    input  [31:0]       reg32_arr__data_in[8],
    output [31:0]       reg32_arr__data_r [8],
    
    // Ports for 'reg16'
    input  [15:0]       reg16__data_in,
    output [15:0]       reg16__data_r ,
    
    // Ports for 'reg8'
    input  [7:0]        reg8__data_in,
    output [7:0]        reg8__data_r 
    
);


// Internal signals
srdl2sv_widget_if #(.ADDR_W (32), .DATA_W(32)) widget_if;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - widget_if -> SystemVerilog interface to between widgets
 *                   and the internal srdl2sv registers.
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA,

     // Interface to internal logic
     .widget_if);

genvar gv_a;


/*******************************************************************
/*******************************************************************
/* REGISTER              : reg32
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        reg32_active     ;
logic        reg32_sw_wr      ;
logic [31:0] reg32_data_mux_in;
logic        reg32_rdy_mux_in ;
logic        reg32_err_mux_in ;
logic [31:0] reg32__data_q    ;


// Register-activation for 'reg32' 
assign reg32_active = widget_if.addr == 0;
assign reg32_sw_wr = reg32_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : data (reg32[31:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge rst_async_n)
if (!rst_async_n)
begin
    reg32__data_q <= 32'd0;
end
else
begin
    if (reg32_sw_wr)
    begin
        if (widget_if.byte_en[0])
            reg32__data_q[7:0] <= widget_if.w_data[7:0];
        if (widget_if.byte_en[1])
            reg32__data_q[15:8] <= widget_if.w_data[15:8];
        if (widget_if.byte_en[2])
            reg32__data_q[23:16] <= widget_if.w_data[23:16];
        if (widget_if.byte_en[3])
            reg32__data_q[31:24] <= widget_if.w_data[31:24];
    end
    else
        // we or wel property not set
        reg32__data_q <= reg32__data_in;
end // of reg32__data's always_ff

// Connect register to hardware output port
assign reg32__data_r = reg32__data_q;




/********************************************** 
 * Assign all fields to signal to Mux         *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg32_data_mux_in = {reg32__data_q};

// Internal registers are ready immediately
assign reg32_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg32_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[3:0])) || (widget_if.w_vld && (|widget_if.byte_en[3:0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg32_arr
/* DIMENSION             : 1
/* DEPTHS (per dimension): [8]
/*******************************************************************
/*******************************************************************/

logic        reg32_arr_active     [8];
logic        reg32_arr_sw_wr      [8];
logic [31:0] reg32_arr_data_mux_in[8];
logic        reg32_arr_rdy_mux_in [8];
logic        reg32_arr_err_mux_in [8];
logic [31:0] reg32_arr__data_q    [8];

generate
for (gv_a = 0; gv_a < 8; gv_a++)
begin
    
    // Register-activation for 'reg32_arr' 
    assign reg32_arr_active[gv_a] = widget_if.addr == 4+(gv_a*4);
    assign reg32_arr_sw_wr[gv_a] = reg32_arr_active[gv_a] && widget_if.w_vld;
    
    //-----------------FIELD SUMMARY-----------------
    // name         : data (reg32_arr[31:0])
    // access       : hw = rw  
    //                sw = rw (precedence)
    // reset        : active_low / asynchronous
    // flags        : ['sw']
    // external     : False
    // storage type : StorageType.FLOPS
    //-----------------------------------------------
    
    always_ff @(posedge clk or negedge rst_async_n)
    if (!rst_async_n)
    begin
        reg32_arr__data_q[gv_a] <= 32'd0;
    end
    else
    begin
        if (reg32_arr_sw_wr[gv_a])
        begin
            if (widget_if.byte_en[0])
                reg32_arr__data_q[gv_a][7:0] <= widget_if.w_data[7:0];
            if (widget_if.byte_en[1])
                reg32_arr__data_q[gv_a][15:8] <= widget_if.w_data[15:8];
            if (widget_if.byte_en[2])
                reg32_arr__data_q[gv_a][23:16] <= widget_if.w_data[23:16];
            if (widget_if.byte_en[3])
                reg32_arr__data_q[gv_a][31:24] <= widget_if.w_data[31:24];
        end
        else
            // we or wel property not set
            reg32_arr__data_q[gv_a] <= reg32_arr__data_in[gv_a];
    end // of reg32_arr__data's always_ff
    
    // Connect register to hardware output port
    assign reg32_arr__data_r[gv_a] = reg32_arr__data_q[gv_a];
    
    
    
    
    /********************************************** 
     * Assign all fields to signal to Mux         *
     **********************************************/
    // Assign all fields. Fields that are not readable are tied to 0.
    assign reg32_arr_data_mux_in[gv_a] = {reg32_arr__data_q[gv_a]};
    
    // Internal registers are ready immediately
    assign reg32_arr_rdy_mux_in[gv_a] = 1'b1;
    
    // Return an error if *no* read and *no* write was succesful. If some bits
    // cannot be read/written but others are succesful, don't return and error
    // Hence, as long as one action can be succesful, no error will be returned.
    assign reg32_arr_err_mux_in[gv_a] = !((widget_if.r_vld && (|widget_if.byte_en[3:0])) || (widget_if.w_vld && (|widget_if.byte_en[3:0])));
end // of for loop with iterator gv_a

endgenerate


/*******************************************************************
/*******************************************************************
/* REGISTER              : reg16
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        reg16_active     ;
logic        reg16_sw_wr      ;
logic [31:0] reg16_data_mux_in;
logic        reg16_rdy_mux_in ;
logic        reg16_err_mux_in ;
logic [15:0] reg16__data_q    ;


// Register-activation for 'reg16' 
assign reg16_active = widget_if.addr == 36;
assign reg16_sw_wr = reg16_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : data (reg16[15:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge rst_async_n)
if (!rst_async_n)
begin
    reg16__data_q <= 16'd0;
end
else
begin
    if (reg16_sw_wr)
    begin
        if (widget_if.byte_en[0])
            reg16__data_q[7:0] <= widget_if.w_data[7:0];
        if (widget_if.byte_en[1])
            reg16__data_q[15:8] <= widget_if.w_data[15:8];
    end
    else
        // we or wel property not set
        reg16__data_q <= reg16__data_in;
end // of reg16__data's always_ff

// Connect register to hardware output port
assign reg16__data_r = reg16__data_q;




/********************************************** 
 * Assign all fields to signal to Mux         *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg16_data_mux_in = {{16{1'b0}}, reg16__data_q};

// Internal registers are ready immediately
assign reg16_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg16_err_mux_in = !((widget_if.r_vld && (|widget_if.byte_en[1:0])) || (widget_if.w_vld && (|widget_if.byte_en[1:0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg8
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        reg8_active     ;
logic [31:0] reg8_data_mux_in;
logic        reg8_rdy_mux_in ;
logic        reg8_err_mux_in ;
logic [7:0]  reg8__data_q    ;


// Register-activation for 'reg8' 
assign reg8_active = widget_if.addr == 40;

//-----------------FIELD SUMMARY-----------------
// name         : data (reg8[7:0])
// access       : hw = rw  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge rst_async_n)
if (!rst_async_n)
begin
    reg8__data_q <= 8'd0;
end
else
begin
        // we or wel property not set
        reg8__data_q <= reg8__data_in;
end // of reg8__data's always_ff

// Connect register to hardware output port
assign reg8__data_r = reg8__data_q;




/********************************************** 
 * Assign all fields to signal to Mux         *
 **********************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg8_data_mux_in = {{24{1'b0}}, reg8__data_q};

// Internal registers are ready immediately
assign reg8_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg8_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (1'b0)));

// Read multiplexer
always_comb
begin
    unique case (1'b1)
        reg32_active:
        begin
            widget_if.r_data = reg32_data_mux_in;
            widget_if.err    = reg32_err_mux_in;
            widget_if.rdy    = reg32_rdy_mux_in;
        end
        reg32_arr_active[0]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[0];
            widget_if.err    = reg32_arr_err_mux_in[0];
            widget_if.rdy    = reg32_arr_rdy_mux_in[0];
        end
        reg32_arr_active[1]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[1];
            widget_if.err    = reg32_arr_err_mux_in[1];
            widget_if.rdy    = reg32_arr_rdy_mux_in[1];
        end
        reg32_arr_active[2]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[2];
            widget_if.err    = reg32_arr_err_mux_in[2];
            widget_if.rdy    = reg32_arr_rdy_mux_in[2];
        end
        reg32_arr_active[3]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[3];
            widget_if.err    = reg32_arr_err_mux_in[3];
            widget_if.rdy    = reg32_arr_rdy_mux_in[3];
        end
        reg32_arr_active[4]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[4];
            widget_if.err    = reg32_arr_err_mux_in[4];
            widget_if.rdy    = reg32_arr_rdy_mux_in[4];
        end
        reg32_arr_active[5]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[5];
            widget_if.err    = reg32_arr_err_mux_in[5];
            widget_if.rdy    = reg32_arr_rdy_mux_in[5];
        end
        reg32_arr_active[6]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[6];
            widget_if.err    = reg32_arr_err_mux_in[6];
            widget_if.rdy    = reg32_arr_rdy_mux_in[6];
        end
        reg32_arr_active[7]:
        begin
            widget_if.r_data = reg32_arr_data_mux_in[7];
            widget_if.err    = reg32_arr_err_mux_in[7];
            widget_if.rdy    = reg32_arr_rdy_mux_in[7];
        end
        reg16_active:
        begin
            widget_if.r_data = reg16_data_mux_in;
            widget_if.err    = reg16_err_mux_in;
            widget_if.rdy    = reg16_rdy_mux_in;
        end
        reg8_active:
        begin
            widget_if.r_data = reg8_data_mux_in;
            widget_if.err    = reg8_err_mux_in;
            widget_if.rdy    = reg8_rdy_mux_in;
        end
        default:
        begin
            // If the address is not found, return an error
            widget_if.r_data = 0;
            widget_if.err    = 1;
            widget_if.rdy    = widget_if.r_vld || widget_if.w_vld;
        end
    endcase
end
endmodule
