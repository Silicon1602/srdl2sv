/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://github.com/Silicon1602/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : October 30 2021 23:34:40
 *  - Path     : /home/dpotter/srdl2sv/examples/hierarchical_regfiles
 *  - RDL file : ['hierarchical_regfiles.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : ./srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : NONE
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Register Bus Type: amba3ahblite
 *  - Address width    : 32
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': False, 'RegFile': False, 'Memory': False, 'Register': False, 'Field': False}
 *
 * ===LICENSE OF HIERARCHICAL_REGFILES.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module hierarchical_regfiles
    
(
    // Resets
     
    
    // Inputs
    input               clk                               ,
    input               HRESETn                           ,
    input  [31:0]       HADDR                             ,
    input               HWRITE                            ,
    input  [2:0]        HSIZE                             ,
    input  [3:0]        HPROT                             ,
    input  [1:0]        HTRANS                            ,
    input  [32-1:0]     HWDATA                            ,
    input               HSEL                              ,
    input  logic        regfile_1__reg_a__f1_hw_wr        ,
    input  logic [15:0] regfile_1__reg_a__f1_in           ,
    input  logic        regfile_1__reg_a__f2_hw_wr        ,
    input  logic [15:0] regfile_1__reg_a__f2_in           ,
    input  logic        regfile_1__reg_b__f1_hw_wr        ,
    input  logic [15:0] regfile_1__reg_b__f1_in           ,
    input  logic        regfile_1__reg_b__f2_hw_wr        ,
    input  logic [15:0] regfile_1__reg_b__f2_in           ,
    input  logic [15:0] regfile_2__regfile_3__reg_d__f1_in[2][4][2],
    input  logic [15:0] regfile_2__regfile_3__reg_d__f2_in[2][4][2],
    input  logic [7:0]  regfile_2__reg_c__f1_in           [2],
    input  logic [15:0] regfile_2__reg_c__f3_in           [2],
    input  logic        reg_e__f1_hw_wr                   ,
    input  logic [15:0] reg_e__f1_in                      ,
    input  logic        reg_e__f2_hw_wr                   ,
    input  logic [15:0] reg_e__f2_in                      ,
    
    // Outputs
    output              HREADYOUT                        ,
    output              HRESP                            ,
    output [32-1:0]     HRDATA                           ,
    output logic [15:0] regfile_1__reg_a__f1_r           ,
    output logic [15:0] regfile_1__reg_a__f2_r           ,
    output logic [15:0] regfile_1__reg_b__f1_r           ,
    output logic [15:0] regfile_1__reg_b__f2_r           ,
    output logic [15:0] regfile_2__regfile_3__reg_d__f1_r[2][4][2],
    output logic [15:0] regfile_2__regfile_3__reg_d__f2_r[2][4][2],
    output logic [7:0]  regfile_2__reg_c__f2_r           [2],
    output logic [15:0] reg_e__f1_r                      ,
    output logic [15:0] reg_e__f2_r                      
);


// Internal signals
srdl2sv_widget_if #(.ADDR_W (32), .DATA_W(32)) widget_if;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - widget_if -> SystemVerilog interface to between widgets
 *                   and the internal srdl2sv registers.
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA,

     // Interface to internal logic
     .widget_if);

genvar gv_a, gv_b, gv_c;

/*******************************************************************
 *******************************************************************
 * REGFILE               : regfile_1
 * DIMENSION             : 0
 * DEPTHS (per dimension): []
 *******************************************************************
 *******************************************************************/


/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_a
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        regfile_1__reg_a_active     ;
logic        regfile_1__reg_a_sw_wr      ;
logic [31:0] regfile_1__reg_a_data_mux_in;
logic        regfile_1__reg_a_rdy_mux_in ;
logic        regfile_1__reg_a_err_mux_in ;
logic [15:0] regfile_1__reg_a__f1_q      ;
logic [15:0] regfile_1__reg_a__f2_q      ;


// Register-activation for 'regfile_1__reg_a' 
assign regfile_1__reg_a_active = widget_if.addr == 0;
assign regfile_1__reg_a_sw_wr = regfile_1__reg_a_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (regfile_1__reg_a[15:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_a_sw_wr)
    begin
        if (widget_if.byte_en[0])
            regfile_1__reg_a__f1_q[7:0] <= widget_if.w_data[7:0];
        if (widget_if.byte_en[1])
            regfile_1__reg_a__f1_q[15:8] <= widget_if.w_data[15:8];
    end
    else
    if (regfile_1__reg_a__f1_hw_wr)
        regfile_1__reg_a__f1_q <= regfile_1__reg_a__f1_in;
end // of regfile_1__reg_a__f1's always_ff

// Connect register to hardware output port
assign regfile_1__reg_a__f1_r = regfile_1__reg_a__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (regfile_1__reg_a[31:16])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_a_sw_wr)
    begin
        if (widget_if.byte_en[2])
            regfile_1__reg_a__f2_q[7:0] <= widget_if.w_data[23:16];
        if (widget_if.byte_en[3])
            regfile_1__reg_a__f2_q[15:8] <= widget_if.w_data[31:24];
    end
    else
    if (regfile_1__reg_a__f2_hw_wr)
        regfile_1__reg_a__f2_q <= regfile_1__reg_a__f2_in;
end // of regfile_1__reg_a__f2's always_ff

// Connect register to hardware output port
assign regfile_1__reg_a__f2_r = regfile_1__reg_a__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign regfile_1__reg_a_data_mux_in = {regfile_1__reg_a__f2_q, regfile_1__reg_a__f1_q};

// Internal registers are ready immediately
assign regfile_1__reg_a_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign regfile_1__reg_a_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])) || (widget_if.w_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_b
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        regfile_1__reg_b_active     ;
logic        regfile_1__reg_b_sw_wr      ;
logic [31:0] regfile_1__reg_b_data_mux_in;
logic        regfile_1__reg_b_rdy_mux_in ;
logic        regfile_1__reg_b_err_mux_in ;
logic [15:0] regfile_1__reg_b__f1_q      ;
logic [15:0] regfile_1__reg_b__f2_q      ;


// Register-activation for 'regfile_1__reg_b' 
assign regfile_1__reg_b_active = widget_if.addr == 4;
assign regfile_1__reg_b_sw_wr = regfile_1__reg_b_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (regfile_1__reg_b[15:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_b_sw_wr)
    begin
        if (widget_if.byte_en[0])
            regfile_1__reg_b__f1_q[7:0] <= widget_if.w_data[7:0];
        if (widget_if.byte_en[1])
            regfile_1__reg_b__f1_q[15:8] <= widget_if.w_data[15:8];
    end
    else
    if (regfile_1__reg_b__f1_hw_wr)
        regfile_1__reg_b__f1_q <= regfile_1__reg_b__f1_in;
end // of regfile_1__reg_b__f1's always_ff

// Connect register to hardware output port
assign regfile_1__reg_b__f1_r = regfile_1__reg_b__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (regfile_1__reg_b[31:16])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (regfile_1__reg_b_sw_wr)
    begin
        if (widget_if.byte_en[2])
            regfile_1__reg_b__f2_q[7:0] <= widget_if.w_data[23:16];
        if (widget_if.byte_en[3])
            regfile_1__reg_b__f2_q[15:8] <= widget_if.w_data[31:24];
    end
    else
    if (regfile_1__reg_b__f2_hw_wr)
        regfile_1__reg_b__f2_q <= regfile_1__reg_b__f2_in;
end // of regfile_1__reg_b__f2's always_ff

// Connect register to hardware output port
assign regfile_1__reg_b__f2_r = regfile_1__reg_b__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign regfile_1__reg_b_data_mux_in = {regfile_1__reg_b__f2_q, regfile_1__reg_b__f1_q};

// Internal registers are ready immediately
assign regfile_1__reg_b_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign regfile_1__reg_b_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])) || (widget_if.w_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])));
/*******************************************************************
 *******************************************************************
 * REGFILE               : regfile_2
 * DIMENSION             : 1
 * DEPTHS (per dimension): [2]
 *******************************************************************
 *******************************************************************/


// Variables of register 'reg_d'
logic        regfile_2__regfile_3__reg_d_active     [2][4][2];
logic        regfile_2__regfile_3__reg_d_sw_wr      [2][4][2];
logic [31:0] regfile_2__regfile_3__reg_d_data_mux_in[2][4][2];
logic        regfile_2__regfile_3__reg_d_rdy_mux_in [2][4][2];
logic        regfile_2__regfile_3__reg_d_err_mux_in [2][4][2];
logic [15:0] regfile_2__regfile_3__reg_d__f1_q      [2][4][2];
logic [15:0] regfile_2__regfile_3__reg_d__f2_q      [2][4][2];

// Variables of register 'reg_c'
logic        regfile_2__reg_c_active     [2];
logic        regfile_2__reg_c_sw_wr      [2];
logic [31:0] regfile_2__reg_c_data_mux_in[2];
logic        regfile_2__reg_c_rdy_mux_in [2];
logic        regfile_2__reg_c_err_mux_in [2];
logic [7:0]  regfile_2__reg_c__f1_q      [2];
logic [7:0]  regfile_2__reg_c__f2_q      [2];
logic [15:0] regfile_2__reg_c__f3_q      [2];

generate
for (gv_a = 0; gv_a < 2; gv_a++)
begin
    /*******************************************************************
     *******************************************************************
     * REGFILE               : regfile_3
     * DIMENSION             : 2
     * DEPTHS (per dimension): [4][2]
     *******************************************************************
     *******************************************************************/
    
    for (gv_b = 0; gv_b < 4; gv_b++)
    begin
        for (gv_c = 0; gv_c < 2; gv_c++)
        begin
            
            /*******************************************************************
            /*******************************************************************
            /* REGISTER              : reg_d
            /* DIMENSION             : 0
            /* DEPTHS (per dimension): []
            /*******************************************************************
            /*******************************************************************/
            
            
            // Register-activation for 'regfile_2__regfile_3__reg_d' 
            assign regfile_2__regfile_3__reg_d_active[gv_a][gv_b][gv_c] = widget_if.addr == 68+(gv_a*36+gv_b*8+gv_c*4);
            assign regfile_2__regfile_3__reg_d_sw_wr[gv_a][gv_b][gv_c] = regfile_2__regfile_3__reg_d_active[gv_a][gv_b][gv_c] && widget_if.w_vld;
            
            //-----------------FIELD SUMMARY-----------------
            // name         : f1 (regfile_2__regfile_3__reg_d[15:0])
            // access       : hw = rw  
            //                sw = rw (precedence)
            // reset        : - / -
            // flags        : ['sw']
            // external     : False
            // storage type : StorageType.FLOPS
            //-----------------------------------------------
            
            always_ff @(posedge clk)
            begin
                if (regfile_2__regfile_3__reg_d_sw_wr[gv_a][gv_b][gv_c])
                begin
                    if (widget_if.byte_en[0])
                        regfile_2__regfile_3__reg_d__f1_q[gv_a][gv_b][gv_c][7:0] <= widget_if.w_data[7:0];
                    if (widget_if.byte_en[1])
                        regfile_2__regfile_3__reg_d__f1_q[gv_a][gv_b][gv_c][15:8] <= widget_if.w_data[15:8];
                end
                else
                    // we or wel property not set
                    regfile_2__regfile_3__reg_d__f1_q[gv_a][gv_b][gv_c] <= regfile_2__regfile_3__reg_d__f1_in[gv_a][gv_b][gv_c];
            end // of regfile_2__regfile_3__reg_d__f1's always_ff
            
            // Connect register to hardware output port
            assign regfile_2__regfile_3__reg_d__f1_r[gv_a][gv_b][gv_c] = regfile_2__regfile_3__reg_d__f1_q[gv_a][gv_b][gv_c];
            
            
            
            //-----------------FIELD SUMMARY-----------------
            // name         : f2 (regfile_2__regfile_3__reg_d[31:16])
            // access       : hw = rw  
            //                sw = rw (precedence)
            // reset        : - / -
            // flags        : ['sw']
            // external     : False
            // storage type : StorageType.FLOPS
            //-----------------------------------------------
            
            always_ff @(posedge clk)
            begin
                if (regfile_2__regfile_3__reg_d_sw_wr[gv_a][gv_b][gv_c])
                begin
                    if (widget_if.byte_en[2])
                        regfile_2__regfile_3__reg_d__f2_q[gv_a][gv_b][gv_c][7:0] <= widget_if.w_data[23:16];
                    if (widget_if.byte_en[3])
                        regfile_2__regfile_3__reg_d__f2_q[gv_a][gv_b][gv_c][15:8] <= widget_if.w_data[31:24];
                end
                else
                    // we or wel property not set
                    regfile_2__regfile_3__reg_d__f2_q[gv_a][gv_b][gv_c] <= regfile_2__regfile_3__reg_d__f2_in[gv_a][gv_b][gv_c];
            end // of regfile_2__regfile_3__reg_d__f2's always_ff
            
            // Connect register to hardware output port
            assign regfile_2__regfile_3__reg_d__f2_r[gv_a][gv_b][gv_c] = regfile_2__regfile_3__reg_d__f2_q[gv_a][gv_b][gv_c];
            
            
            
            
            /************************************** 
             * Assign all fields to signal to Mux *
             **************************************/
            // Assign all fields. Fields that are not readable are tied to 0.
            assign regfile_2__regfile_3__reg_d_data_mux_in[gv_a][gv_b][gv_c] = {regfile_2__regfile_3__reg_d__f2_q[gv_a][gv_b][gv_c], regfile_2__regfile_3__reg_d__f1_q[gv_a][gv_b][gv_c]};
            
            // Internal registers are ready immediately
            assign regfile_2__regfile_3__reg_d_rdy_mux_in[gv_a][gv_b][gv_c] = 1'b1;
            
            // Return an error if *no* read and *no* write was succesful. If some bits
            // cannot be read/written but others are succesful, don't return and error
            // Hence, as long as one action can be succesful, no error will be returned.
            assign regfile_2__regfile_3__reg_d_err_mux_in[gv_a][gv_b][gv_c] = !((widget_if.r_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])) || (widget_if.w_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])));
        end // of for loop with iterator gv_b
    end // of for loop with iterator gv_a
    
    /*******************************************************************
    /*******************************************************************
    /* REGISTER              : reg_c
    /* DIMENSION             : 0
    /* DEPTHS (per dimension): []
    /*******************************************************************
    /*******************************************************************/
    
    
    // Register-activation for 'regfile_2__reg_c' 
    assign regfile_2__reg_c_active[gv_a] = widget_if.addr == 64+(gv_a*36);
    assign regfile_2__reg_c_sw_wr[gv_a] = regfile_2__reg_c_active[gv_a] && widget_if.w_vld;
    
    //-----------------FIELD SUMMARY-----------------
    // name         : f1 (regfile_2__reg_c[7:0])
    // access       : hw = w  
    //                sw = r (precedence)
    // reset        : - / -
    // flags        : ['sw']
    // external     : False
    // storage type : StorageType.WIRE
    //-----------------------------------------------
    
    // Field is a simple wire.
    // To generate a flop either add the we/wel property, add
    // a reset, or change the sw/hw access properties
    assign regfile_2__reg_c__f1_q[gv_a] = regfile_2__reg_c__f1_in[gv_a];
    
    //-----------------FIELD SUMMARY-----------------
    // name         : f2 (regfile_2__reg_c[15:8])
    // access       : hw = r  
    //                sw = r (precedence)
    // reset        : - / -
    // flags        : ['sw']
    // external     : False
    // storage type : StorageType.CONST
    //-----------------------------------------------
    
    // Field is defined as a constant.
    assign regfile_2__reg_c__f2_q[gv_a] = 8'd42;
    
    // Connect register to hardware output port
    assign regfile_2__reg_c__f2_r[gv_a] = regfile_2__reg_c__f2_q[gv_a];
    
    //-----------------FIELD SUMMARY-----------------
    // name         : f3 (regfile_2__reg_c[31:16])
    // access       : hw = w  
    //                sw = rw (precedence)
    // reset        : - / -
    // flags        : ['sw']
    // external     : False
    // storage type : StorageType.FLOPS
    //-----------------------------------------------
    
    always_ff @(posedge clk)
    begin
        if (regfile_2__reg_c_sw_wr[gv_a])
        begin
            if (widget_if.byte_en[2])
                regfile_2__reg_c__f3_q[gv_a][7:0] <= widget_if.w_data[23:16];
            if (widget_if.byte_en[3])
                regfile_2__reg_c__f3_q[gv_a][15:8] <= widget_if.w_data[31:24];
        end
        else
            // we or wel property not set
            regfile_2__reg_c__f3_q[gv_a] <= regfile_2__reg_c__f3_in[gv_a];
    end // of regfile_2__reg_c__f3's always_ff
    
    
    
    
    /************************************** 
     * Assign all fields to signal to Mux *
     **************************************/
    // Assign all fields. Fields that are not readable are tied to 0.
    assign regfile_2__reg_c_data_mux_in[gv_a] = {regfile_2__reg_c__f3_q[gv_a], regfile_2__reg_c__f2_q[gv_a], regfile_2__reg_c__f1_q[gv_a]};
    
    // Internal registers are ready immediately
    assign regfile_2__reg_c_rdy_mux_in[gv_a] = 1'b1;
    
    // Return an error if *no* read and *no* write was succesful. If some bits
    // cannot be read/written but others are succesful, don't return and error
    // Hence, as long as one action can be succesful, no error will be returned.
    assign regfile_2__reg_c_err_mux_in[gv_a] = !((widget_if.r_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])) || (widget_if.w_vld && (widget_if.byte_en[2] || widget_if.byte_en[3])));
end // of for loop with iterator gv_a
endgenerate


/*******************************************************************
/*******************************************************************
/* REGISTER              : reg_e
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        reg_e_active     ;
logic        reg_e_sw_wr      ;
logic [31:0] reg_e_data_mux_in;
logic        reg_e_rdy_mux_in ;
logic        reg_e_err_mux_in ;
logic [15:0] reg_e__f1_q      ;
logic [15:0] reg_e__f2_q      ;


// Register-activation for 'reg_e' 
assign reg_e_active = widget_if.addr == 136;
assign reg_e_sw_wr = reg_e_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : f1 (reg_e[15:0])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_e_sw_wr)
    begin
        if (widget_if.byte_en[0])
            reg_e__f1_q[7:0] <= widget_if.w_data[7:0];
        if (widget_if.byte_en[1])
            reg_e__f1_q[15:8] <= widget_if.w_data[15:8];
    end
    else
    if (reg_e__f1_hw_wr)
        reg_e__f1_q <= reg_e__f1_in;
end // of reg_e__f1's always_ff

// Connect register to hardware output port
assign reg_e__f1_r = reg_e__f1_q;



//-----------------FIELD SUMMARY-----------------
// name         : f2 (reg_e[31:16])
// access       : hw = rw  
//                sw = rw (precedence)
// reset        : - / -
// flags        : ['sw', 'we']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (reg_e_sw_wr)
    begin
        if (widget_if.byte_en[2])
            reg_e__f2_q[7:0] <= widget_if.w_data[23:16];
        if (widget_if.byte_en[3])
            reg_e__f2_q[15:8] <= widget_if.w_data[31:24];
    end
    else
    if (reg_e__f2_hw_wr)
        reg_e__f2_q <= reg_e__f2_in;
end // of reg_e__f2's always_ff

// Connect register to hardware output port
assign reg_e__f2_r = reg_e__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign reg_e_data_mux_in = {reg_e__f2_q, reg_e__f1_q};

// Internal registers are ready immediately
assign reg_e_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign reg_e_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])) || (widget_if.w_vld && (widget_if.byte_en[0] || widget_if.byte_en[1] || widget_if.byte_en[2] || widget_if.byte_en[3])));

// Read multiplexer
always_comb
begin
    unique case (1'b1)
        regfile_1__reg_a_active:
        begin
            widget_if.r_data = regfile_1__reg_a_data_mux_in;
            widget_if.err    = regfile_1__reg_a_err_mux_in;
            widget_if.rdy    = regfile_1__reg_a_rdy_mux_in;
        end
        regfile_1__reg_b_active:
        begin
            widget_if.r_data = regfile_1__reg_b_data_mux_in;
            widget_if.err    = regfile_1__reg_b_err_mux_in;
            widget_if.rdy    = regfile_1__reg_b_rdy_mux_in;
        end
        regfile_2__regfile_3__reg_d_active[0][0][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][0][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][0][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][0][0];
        end
        regfile_2__regfile_3__reg_d_active[0][0][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][0][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][0][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][0][1];
        end
        regfile_2__regfile_3__reg_d_active[0][1][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][1][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][1][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][1][0];
        end
        regfile_2__regfile_3__reg_d_active[0][1][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][1][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][1][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][1][1];
        end
        regfile_2__regfile_3__reg_d_active[0][2][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][2][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][2][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][2][0];
        end
        regfile_2__regfile_3__reg_d_active[0][2][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][2][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][2][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][2][1];
        end
        regfile_2__regfile_3__reg_d_active[0][3][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][3][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][3][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][3][0];
        end
        regfile_2__regfile_3__reg_d_active[0][3][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[0][3][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[0][3][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[0][3][1];
        end
        regfile_2__regfile_3__reg_d_active[1][0][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][0][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][0][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][0][0];
        end
        regfile_2__regfile_3__reg_d_active[1][0][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][0][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][0][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][0][1];
        end
        regfile_2__regfile_3__reg_d_active[1][1][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][1][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][1][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][1][0];
        end
        regfile_2__regfile_3__reg_d_active[1][1][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][1][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][1][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][1][1];
        end
        regfile_2__regfile_3__reg_d_active[1][2][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][2][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][2][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][2][0];
        end
        regfile_2__regfile_3__reg_d_active[1][2][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][2][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][2][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][2][1];
        end
        regfile_2__regfile_3__reg_d_active[1][3][0]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][3][0];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][3][0];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][3][0];
        end
        regfile_2__regfile_3__reg_d_active[1][3][1]:
        begin
            widget_if.r_data = regfile_2__regfile_3__reg_d_data_mux_in[1][3][1];
            widget_if.err    = regfile_2__regfile_3__reg_d_err_mux_in[1][3][1];
            widget_if.rdy    = regfile_2__regfile_3__reg_d_rdy_mux_in[1][3][1];
        end
        regfile_2__reg_c_active[0]:
        begin
            widget_if.r_data = regfile_2__reg_c_data_mux_in[0];
            widget_if.err    = regfile_2__reg_c_err_mux_in[0];
            widget_if.rdy    = regfile_2__reg_c_rdy_mux_in[0];
        end
        regfile_2__reg_c_active[1]:
        begin
            widget_if.r_data = regfile_2__reg_c_data_mux_in[1];
            widget_if.err    = regfile_2__reg_c_err_mux_in[1];
            widget_if.rdy    = regfile_2__reg_c_rdy_mux_in[1];
        end
        reg_e_active:
        begin
            widget_if.r_data = reg_e_data_mux_in;
            widget_if.err    = reg_e_err_mux_in;
            widget_if.rdy    = reg_e_rdy_mux_in;
        end
        default:
        begin
            // If the address is not found, return an error
            widget_if.r_data = 0;
            widget_if.err    = 1;
            widget_if.rdy    = widget_if.r_vld || widget_if.w_vld;
        end
    endcase
end
endmodule
