package enums_pkg;

typedef enum logic [1:0] {
    val_1 = 2'd2,
    val_2 = 2'd1
} first_enum;

typedef enum logic [1:0] {
    val_3 = 2'd2,
    val_4 = 2'd1
} second_enum;

typedef enum logic [1:0] {
    val_5 = 2'd2,
    val_6 = 2'd1
} third_enum;

endpackage
