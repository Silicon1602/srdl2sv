/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://git.dennispotter.eu/Dennis/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : October 20 2021 23:49:07
 *  - Path     : /home/dpotter/srdl2sv_second_repo/examples/simple_rw_reg
 *  - RDL file : ['simple_rw_reg.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : ./srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : INFO
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Register Bus Type: amba3ahblite
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': False, 'RegFile': False, 'Memory': False, 'Register': False, 'Field': False}
 *
 * ===LICENSE OF SIMPLE_RW_REG.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module simple_rw_reg
    import srdl2sv_if_pkg::*;
(
    // Resets
     
    
    // Inputs
    input               clk                  ,
    input               HRESETn              ,
    input  [31:0]       HADDR                ,
    input               HWRITE               ,
    input  [2:0]        HSIZE                ,
    input  [3:0]        HPROT                ,
    input  [1:0]        HTRANS               ,
    input  [32-1:0]     HWDATA               ,
    input               HSEL                 ,
    input  logic        register_1d__f1_hw_wr,
    input  logic [15:0] register_1d__f1_in   ,
    input  logic        register_1d__f2_hw_wr,
    input  logic [15:0] register_1d__f2_in   ,
    input  logic        register_2d__f1_hw_wr[2],
    input  logic [15:0] register_2d__f1_in   [2],
    input  logic        register_2d__f2_hw_wr[2],
    input  logic [15:0] register_2d__f2_in   [2],
    input  logic        register_3d__f1_hw_wr[2][2],
    input  logic [15:0] register_3d__f1_in   [2][2],
    input  logic        register_3d__f2_hw_wr[2][2],
    input  logic [15:0] register_3d__f2_in   [2][2],
    
    // Outputs
    output              HREADYOUT        ,
    output              HRESP            ,
    output [32-1:0]     HRDATA           ,
    output logic [15:0] register_1d__f1_r,
    output logic [15:0] register_1d__f2_r,
    output logic [15:0] register_2d__f1_r[2],
    output logic [15:0] register_2d__f2_r[2],
    output logic [15:0] register_3d__f1_r[2][2],
    output logic [15:0] register_3d__f2_r[2][2]
);


// Internal signals
b2r_t b2r;
r2b_t r2b;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - r2b.*     -> Signals from registers to bus
 *    - b2r.*     -> Signals from bus to registers
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Outputs to internal logic
     .b2r,

     // Inputs from internal logic
     .r2b,

     // Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA);

genvar gv_a, gv_b;


/*******************************************************************
/*******************************************************************
/* REGISTER              : register_1d
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        register_1d_active     ;
logic        register_1d_sw_wr      ;
logic [31:0] register_1d_data_mux_in;
logic        register_1d_rdy_mux_in ;
logic        register_1d_err_mux_in ;
logic [15:0] register_1d__f1_q      ;
logic [15:0] register_1d__f2_q      ;


// Register-activation for 'register_1d' 
assign register_1d_active = b2r.addr == 0;
assign register_1d_sw_wr = register_1d_active && b2r.w_vld;

//-----------------FIELD SUMMARY-----------------
// name       : f1 (register_1d[15:0])
// access     : hw = rw  
//              sw = rw (precedence)
// reset      : - / -
// flags      : ['sw', 'we']
// external   : False
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (register_1d_sw_wr)
    begin
        if (b2r.byte_en[0])
            register_1d__f1_q[7:0] <= b2r.data[7:0];
        if (b2r.byte_en[1])
            register_1d__f1_q[15:8] <= b2r.data[15:8];
    end
    else
    if (register_1d__f1_hw_wr)
        register_1d__f1_q <= register_1d__f1_in;
end // of register_1d__f1's always_ff

// Connect register to hardware output port
assign register_1d__f1_r = register_1d__f1_q;



//-----------------FIELD SUMMARY-----------------
// name       : f2 (register_1d[31:16])
// access     : hw = rw  
//              sw = rw (precedence)
// reset      : - / -
// flags      : ['sw', 'we']
// external   : False
//-----------------------------------------------

always_ff @(posedge clk)
begin
    if (register_1d_sw_wr)
    begin
        if (b2r.byte_en[2])
            register_1d__f2_q[7:0] <= b2r.data[23:16];
        if (b2r.byte_en[3])
            register_1d__f2_q[15:8] <= b2r.data[31:24];
    end
    else
    if (register_1d__f2_hw_wr)
        register_1d__f2_q <= register_1d__f2_in;
end // of register_1d__f2's always_ff

// Connect register to hardware output port
assign register_1d__f2_r = register_1d__f2_q;




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign register_1d_data_mux_in = {register_1d__f2_q, register_1d__f1_q};

// Internal registers are ready immediately
assign register_1d_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign register_1d_err_mux_in = !((b2r.r_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])) || (b2r.w_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : register_2d
/* DIMENSION             : 1
/* DEPTHS (per dimension): [2]
/*******************************************************************
/*******************************************************************/

logic        register_2d_active     [2];
logic        register_2d_sw_wr      [2];
logic [31:0] register_2d_data_mux_in[2];
logic        register_2d_rdy_mux_in [2];
logic        register_2d_err_mux_in [2];
logic [15:0] register_2d__f1_q      [2];
logic [15:0] register_2d__f2_q      [2];

generate
for (gv_a = 0; gv_a < 2; gv_a++)
begin
    
    // Register-activation for 'register_2d' 
    assign register_2d_active[gv_a] = b2r.addr == 4+(gv_a*4);
    assign register_2d_sw_wr[gv_a] = register_2d_active[gv_a] && b2r.w_vld;
    
    //-----------------FIELD SUMMARY-----------------
    // name       : f1 (register_2d[15:0])
    // access     : hw = rw  
    //              sw = rw (precedence)
    // reset      : - / -
    // flags      : ['sw', 'we']
    // external   : False
    //-----------------------------------------------
    
    always_ff @(posedge clk)
    begin
        if (register_2d_sw_wr[gv_a])
        begin
            if (b2r.byte_en[0])
                register_2d__f1_q[gv_a][7:0] <= b2r.data[7:0];
            if (b2r.byte_en[1])
                register_2d__f1_q[gv_a][15:8] <= b2r.data[15:8];
        end
        else
        if (register_2d__f1_hw_wr[gv_a])
            register_2d__f1_q[gv_a] <= register_2d__f1_in[gv_a];
    end // of register_2d__f1's always_ff
    
    // Connect register to hardware output port
    assign register_2d__f1_r[gv_a] = register_2d__f1_q[gv_a];
    
    
    
    //-----------------FIELD SUMMARY-----------------
    // name       : f2 (register_2d[31:16])
    // access     : hw = rw  
    //              sw = rw (precedence)
    // reset      : - / -
    // flags      : ['sw', 'we']
    // external   : False
    //-----------------------------------------------
    
    always_ff @(posedge clk)
    begin
        if (register_2d_sw_wr[gv_a])
        begin
            if (b2r.byte_en[2])
                register_2d__f2_q[gv_a][7:0] <= b2r.data[23:16];
            if (b2r.byte_en[3])
                register_2d__f2_q[gv_a][15:8] <= b2r.data[31:24];
        end
        else
        if (register_2d__f2_hw_wr[gv_a])
            register_2d__f2_q[gv_a] <= register_2d__f2_in[gv_a];
    end // of register_2d__f2's always_ff
    
    // Connect register to hardware output port
    assign register_2d__f2_r[gv_a] = register_2d__f2_q[gv_a];
    
    
    
    
    /************************************** 
     * Assign all fields to signal to Mux *
     **************************************/
    // Assign all fields. Fields that are not readable are tied to 0.
    assign register_2d_data_mux_in[gv_a] = {register_2d__f2_q[gv_a], register_2d__f1_q[gv_a]};
    
    // Internal registers are ready immediately
    assign register_2d_rdy_mux_in[gv_a] = 1'b1;
    
    // Return an error if *no* read and *no* write was succesful. If some bits
    // cannot be read/written but others are succesful, don't return and error
    // Hence, as long as one action can be succesful, no error will be returned.
    assign register_2d_err_mux_in[gv_a] = !((b2r.r_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])) || (b2r.w_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])));
end // of for loop with iterator gv_a

endgenerate


/*******************************************************************
/*******************************************************************
/* REGISTER              : register_3d
/* DIMENSION             : 2
/* DEPTHS (per dimension): [2][2]
/*******************************************************************
/*******************************************************************/

logic        register_3d_active     [2][2];
logic        register_3d_sw_wr      [2][2];
logic [31:0] register_3d_data_mux_in[2][2];
logic        register_3d_rdy_mux_in [2][2];
logic        register_3d_err_mux_in [2][2];
logic [15:0] register_3d__f1_q      [2][2];
logic [15:0] register_3d__f2_q      [2][2];

generate
for (gv_a = 0; gv_a < 2; gv_a++)
begin
    for (gv_b = 0; gv_b < 2; gv_b++)
    begin
        
        // Register-activation for 'register_3d' 
        assign register_3d_active[gv_a][gv_b] = b2r.addr == 12+(gv_a*8+gv_b*4);
        assign register_3d_sw_wr[gv_a][gv_b] = register_3d_active[gv_a][gv_b] && b2r.w_vld;
        
        //-----------------FIELD SUMMARY-----------------
        // name       : f1 (register_3d[15:0])
        // access     : hw = rw  
        //              sw = rw (precedence)
        // reset      : - / -
        // flags      : ['sw', 'we']
        // external   : False
        //-----------------------------------------------
        
        always_ff @(posedge clk)
        begin
            if (register_3d_sw_wr[gv_a][gv_b])
            begin
                if (b2r.byte_en[0])
                    register_3d__f1_q[gv_a][gv_b][7:0] <= b2r.data[7:0];
                if (b2r.byte_en[1])
                    register_3d__f1_q[gv_a][gv_b][15:8] <= b2r.data[15:8];
            end
            else
            if (register_3d__f1_hw_wr[gv_a][gv_b])
                register_3d__f1_q[gv_a][gv_b] <= register_3d__f1_in[gv_a][gv_b];
        end // of register_3d__f1's always_ff
        
        // Connect register to hardware output port
        assign register_3d__f1_r[gv_a][gv_b] = register_3d__f1_q[gv_a][gv_b];
        
        
        
        //-----------------FIELD SUMMARY-----------------
        // name       : f2 (register_3d[31:16])
        // access     : hw = rw  
        //              sw = rw (precedence)
        // reset      : - / -
        // flags      : ['sw', 'we']
        // external   : False
        //-----------------------------------------------
        
        always_ff @(posedge clk)
        begin
            if (register_3d_sw_wr[gv_a][gv_b])
            begin
                if (b2r.byte_en[2])
                    register_3d__f2_q[gv_a][gv_b][7:0] <= b2r.data[23:16];
                if (b2r.byte_en[3])
                    register_3d__f2_q[gv_a][gv_b][15:8] <= b2r.data[31:24];
            end
            else
            if (register_3d__f2_hw_wr[gv_a][gv_b])
                register_3d__f2_q[gv_a][gv_b] <= register_3d__f2_in[gv_a][gv_b];
        end // of register_3d__f2's always_ff
        
        // Connect register to hardware output port
        assign register_3d__f2_r[gv_a][gv_b] = register_3d__f2_q[gv_a][gv_b];
        
        
        
        
        /************************************** 
         * Assign all fields to signal to Mux *
         **************************************/
        // Assign all fields. Fields that are not readable are tied to 0.
        assign register_3d_data_mux_in[gv_a][gv_b] = {register_3d__f2_q[gv_a][gv_b], register_3d__f1_q[gv_a][gv_b]};
        
        // Internal registers are ready immediately
        assign register_3d_rdy_mux_in[gv_a][gv_b] = 1'b1;
        
        // Return an error if *no* read and *no* write was succesful. If some bits
        // cannot be read/written but others are succesful, don't return and error
        // Hence, as long as one action can be succesful, no error will be returned.
        assign register_3d_err_mux_in[gv_a][gv_b] = !((b2r.r_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])) || (b2r.w_vld && (b2r.byte_en[0] || b2r.byte_en[1] || b2r.byte_en[2] || b2r.byte_en[3])));
    end // of for loop with iterator gv_b
end // of for loop with iterator gv_a

endgenerate


// Read multiplexer
always_comb
begin
    unique case (1'b1)
        register_1d_active:
        begin
            r2b.data = register_1d_data_mux_in;
            r2b.err  = register_1d_err_mux_in;
            r2b.rdy  = register_1d_rdy_mux_in;
        end
        register_2d_active[0]:
        begin
            r2b.data = register_2d_data_mux_in[0];
            r2b.err  = register_2d_err_mux_in[0];
            r2b.rdy  = register_2d_rdy_mux_in[0];
        end
        register_2d_active[1]:
        begin
            r2b.data = register_2d_data_mux_in[1];
            r2b.err  = register_2d_err_mux_in[1];
            r2b.rdy  = register_2d_rdy_mux_in[1];
        end
        register_3d_active[0][0]:
        begin
            r2b.data = register_3d_data_mux_in[0][0];
            r2b.err  = register_3d_err_mux_in[0][0];
            r2b.rdy  = register_3d_rdy_mux_in[0][0];
        end
        register_3d_active[0][1]:
        begin
            r2b.data = register_3d_data_mux_in[0][1];
            r2b.err  = register_3d_err_mux_in[0][1];
            r2b.rdy  = register_3d_rdy_mux_in[0][1];
        end
        register_3d_active[1][0]:
        begin
            r2b.data = register_3d_data_mux_in[1][0];
            r2b.err  = register_3d_err_mux_in[1][0];
            r2b.rdy  = register_3d_rdy_mux_in[1][0];
        end
        register_3d_active[1][1]:
        begin
            r2b.data = register_3d_data_mux_in[1][1];
            r2b.err  = register_3d_err_mux_in[1][1];
            r2b.rdy  = register_3d_rdy_mux_in[1][1];
        end
        default:
        begin
            // If the address is not found, return an error
            r2b.data = 0;
            r2b.err  = 1;
            r2b.rdy  = b2r.r_vld || b2r.w_vld;
        end
    endcase
end
endmodule
