package enums__regfile_1_pkg;

typedef enum logic [1:0] {
    val_7 = 2'd2,
    val_8 = 2'd1
} fourth_enum;

endpackage
