module {addrmap_name} (
    {bus_io}
    {io_list}
);

    {bus_widget}

    {registers}
endmodule
