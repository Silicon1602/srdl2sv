/*****************************************************************
 *
 *    ███████╗██████╗ ██████╗ ██╗     ██████╗ ███████╗██╗   ██╗
 *    ██╔════╝██╔══██╗██╔══██╗██║     ╚════██╗██╔════╝██║   ██║
 *    ███████╗██████╔╝██║  ██║██║      █████╔╝███████╗██║   ██║
 *    ╚════██║██╔══██╗██║  ██║██║     ██╔═══╝ ╚════██║╚██╗ ██╔╝
 *    ███████║██║  ██║██████╔╝███████╗███████╗███████║ ╚████╔╝ 
 *    ╚══════╝╚═╝  ╚═╝╚═════╝ ╚══════╝╚══════╝╚══════╝  ╚═══╝  
 *
 * The present RTL was generated by srdl2sv v0.01. The RTL and all
 * templates the RTL is derived from are licensed under the MIT
 * license. The license is shown below.
 *
 * srdl2sv itself is licensed under GPLv3.
 *
 * Maintainer : Dennis Potter <dennis@dennispotter.eu>
 * Report Bugs: https://github.com/Silicon1602/srdl2sv/issues
 *
 * ===GENERATION INFORMATION======================================
 *
 * Generation information:
 *  - User:    : dpotter
 *  - Time     : October 30 2021 23:34:49
 *  - Path     : /home/dpotter/srdl2sv/examples/interrupt_hierarchy
 *  - RDL file : ['interrupt_hierarchy.rdl']
 *  - Hostname : ArchXPS 
 * 
 * RDL include directories:
 *  - 
 *
 * Commandline arguments to srdl2sv:
 *  - Ouput Directory  : ./srdl2sv_out
 *  - Stream Log Level : INFO
 *  - File Log Level   : NONE
 *  - Use Real Tabs    : False
 *  - Tab Width        : 4
 *  - Enums Enabled    : True
 *  - Register Bus Type: amba3ahblite
 *  - Address width    : 32
 *  - Byte enables     : True
 *  - Descriptions     : {'AddrMap': False, 'RegFile': False, 'Memory': False, 'Register': False, 'Field': False}
 *
 * ===LICENSE OF INTERRUPT_HIERARCHY.SV=====================================
 *
 * Copyright 2021 Dennis Potter <dennis@dennispotter.eu>
 * 
 * Permission is hereby granted, free of charge, to any person 
 * obtaining a copy of this software and associated documentation
 * files (the "Software"), to deal in the Software without 
 * restriction, including without limitation the rights to use, 
 * copy, modify, merge, publish, distribute, sublicense, and/or 
 * sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following 
 * conditions:
 * 
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
 * OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
 * NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
 * WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
 * OTHER DEALINGS IN THE SOFTWARE.
 ****************************************************************/
module interrupt_hierarchy
    
(
    // Resets
    input  field_reset_n, 
    
    // Inputs
    input              clk                                ,
    input              HRESETn                            ,
    input  [31:0]      HADDR                              ,
    input              HWRITE                             ,
    input  [2:0]       HSIZE                              ,
    input  [3:0]       HPROT                              ,
    input  [1:0]       HTRANS                             ,
    input  [32-1:0]    HWDATA                             ,
    input              HSEL                               ,
    input  logic [0:0] block_a_int__crc_error_in          ,
    input  logic [0:0] block_a_int__len_error_in          ,
    input  logic [0:0] block_a_int__multi_bit_ecc_error_in,
    input  logic [3:0] block_a_int__active_ecc_master_in  ,
    input  logic [0:0] block_b_int__crc_error_in          ,
    input  logic [0:0] block_b_int__len_error_in          ,
    input  logic [0:0] block_b_int__multi_bit_ecc_error_in,
    input  logic [3:0] block_b_int__active_ecc_master_in  ,
    input  logic [0:0] block_c_int__crc_error_in          ,
    input  logic [0:0] block_c_int__len_error_in          ,
    input  logic [0:0] block_c_int__multi_bit_ecc_error_in,
    input  logic [3:0] block_c_int__active_ecc_master_in  ,
    input  logic [0:0] block_d_int__crc_error_in          ,
    input  logic [0:0] block_d_int__len_error_in          ,
    input  logic [0:0] block_d_int__multi_bit_ecc_error_in,
    input  logic [3:0] block_d_int__active_ecc_master_in  ,
    
    // Outputs
    output          HREADYOUT       ,
    output          HRESP           ,
    output [32-1:0] HRDATA          ,
    output logic    block_a_int_intr,
    output logic    block_a_int_halt,
    output logic    block_b_int_intr,
    output logic    block_b_int_halt,
    output logic    block_c_int_intr,
    output logic    block_c_int_halt,
    output logic    block_d_int_intr,
    output logic    block_d_int_halt,
    output logic    master_int_intr ,
    output logic    master_halt_intr,
    output logic    master_halt_halt,
    output logic    global_int_intr ,
    output logic    global_int_halt 
);


// Internal signals
srdl2sv_widget_if #(.ADDR_W (32), .DATA_W(32)) widget_if;

/*******************************************************************
 * AMBA 3 AHB Lite Widget
 * ======================
 * Naming conventions
 *    - widget_if -> SystemVerilog interface to between widgets
 *                   and the internal srdl2sv registers.
 *    - H*        -> Signals as defined in AMBA3 AHB Lite 
 *                   specification
 *    - clk       -> Clock that drives registers and the bus
 *******************************************************************/
srdl2sv_amba3ahblite
     #(.FLOP_REGISTER_IF (0),
       .BUS_BITS         (32),
       .NO_BYTE_ENABLE   (0))
srdl2sv_amba3ahblite_inst
     (// Bus protocol
     .HRESETn,
     .HCLK        (clk),
     .HADDR,
     .HWRITE,
     .HSIZE,
     .HPROT,
     .HTRANS,
     .HWDATA,
     .HSEL,

     .HREADYOUT,
     .HRESP,
     .HRDATA,

     // Interface to internal logic
     .widget_if);

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_a_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_a_int_active                      ;
logic        block_a_int_sw_wr                       ;
logic [31:0] block_a_int_data_mux_in                 ;
logic        block_a_int_rdy_mux_in                  ;
logic        block_a_int_err_mux_in                  ;
logic [0:0]  block_a_int__crc_error_q                ;
logic [0:0]  block_a_int__crc_error_sticky_latch     ;
logic [0:0]  block_a_int__len_error_q                ;
logic [0:0]  block_a_int__len_error_sticky_latch     ;
logic [0:0]  block_a_int__multi_bit_ecc_error_q      ;
logic [0:0]  block_a_int__multi_bit_ecc_error_sticky_latch;
logic [3:0]  block_a_int__active_ecc_master_q        ;
logic [3:0]  block_a_int__active_ecc_master_sticky_latch;


// Register-activation for 'block_a_int' 
assign block_a_int_active = widget_if.addr == 0;
assign block_a_int_sw_wr = block_a_int_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_a_int[0:0])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int__crc_error_q <= 1'd0;
end
else
begin
    if (block_a_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_a_int__crc_error_q[0:0] <= block_a_int__crc_error_q[0:0] & ~widget_if.w_data[0:0];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_a_int__crc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_a_int__crc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_a_int__crc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_a_int__crc_error_sticky_latch = block_a_int__crc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_a_int[1:1])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int__len_error_q <= 1'd0;
end
else
begin
    if (block_a_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_a_int__len_error_q[0:0] <= block_a_int__len_error_q[0:0] & ~widget_if.w_data[1:1];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_a_int__len_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_a_int__len_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_a_int__len_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_a_int__len_error_sticky_latch = block_a_int__len_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_a_int[2:2])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_a_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_a_int__multi_bit_ecc_error_q[0:0] <= block_a_int__multi_bit_ecc_error_q[0:0] & ~widget_if.w_data[2:2];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_a_int__multi_bit_ecc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_a_int__multi_bit_ecc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_a_int__multi_bit_ecc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_a_int__multi_bit_ecc_error_sticky_latch = block_a_int__multi_bit_ecc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : active_ecc_master (block_a_int[7:4])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'sticky']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int__active_ecc_master_q <= 4'd0;
end
else
begin
    if (block_a_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_a_int__active_ecc_master_q[3:0] <= block_a_int__active_ecc_master_q[3:0] & ~widget_if.w_data[7:4];
        end
    end
    else
    if (|block_a_int__active_ecc_master_sticky_latch && !(|block_a_int__active_ecc_master_q))
    begin
        // Sticky. Keep value until software clears it
        block_a_int__active_ecc_master_q <= block_a_int__active_ecc_master_in;
    end
end // of block_a_int__active_ecc_master's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_a_int__active_ecc_master_sticky_latch = block_a_int__active_ecc_master_in;


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign block_a_int_intr = |(block_a_int__crc_error_q & block_a_int_en__crc_error_q) || |(block_a_int__len_error_q & block_a_int_en__len_error_q) || |(block_a_int__multi_bit_ecc_error_q & block_a_int_en__multi_bit_ecc_error_q);

// Register has at least one interrupt field with halt property set
assign block_a_int_halt = |(block_a_int__crc_error_q & ~block_a_halt_en__crc_error_q) || |(block_a_int__len_error_q & ~block_a_halt_en__len_error_q) || |(block_a_int__multi_bit_ecc_error_q & ~block_a_halt_en__multi_bit_ecc_error_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_a_int_data_mux_in = {{24{1'b0}}, block_a_int__active_ecc_master_q, {1{1'b0}}, block_a_int__multi_bit_ecc_error_q, block_a_int__len_error_q, block_a_int__crc_error_q};

// Internal registers are ready immediately
assign block_a_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_a_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_a_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_a_int_en_active                ;
logic        block_a_int_en_sw_wr                 ;
logic [31:0] block_a_int_en_data_mux_in           ;
logic        block_a_int_en_rdy_mux_in            ;
logic        block_a_int_en_err_mux_in            ;
logic [0:0]  block_a_int_en__crc_error_q          ;
logic [0:0]  block_a_int_en__len_error_q          ;
logic [0:0]  block_a_int_en__multi_bit_ecc_error_q;


// Register-activation for 'block_a_int_en' 
assign block_a_int_en_active = widget_if.addr == 4;
assign block_a_int_en_sw_wr = block_a_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_a_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int_en__crc_error_q <= 1'd1;
end
else
begin
    if (block_a_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_int_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_a_int_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_a_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int_en__len_error_q <= 1'd1;
end
else
begin
    if (block_a_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_int_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_a_int_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_a_int_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_int_en__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_a_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_int_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_a_int_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_a_int_en_data_mux_in = {{29{1'b0}}, block_a_int_en__multi_bit_ecc_error_q, block_a_int_en__len_error_q, block_a_int_en__crc_error_q};

// Internal registers are ready immediately
assign block_a_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_a_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_a_halt_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_a_halt_en_active                ;
logic        block_a_halt_en_sw_wr                 ;
logic [31:0] block_a_halt_en_data_mux_in           ;
logic        block_a_halt_en_rdy_mux_in            ;
logic        block_a_halt_en_err_mux_in            ;
logic [0:0]  block_a_halt_en__crc_error_q          ;
logic [0:0]  block_a_halt_en__len_error_q          ;
logic [0:0]  block_a_halt_en__multi_bit_ecc_error_q;


// Register-activation for 'block_a_halt_en' 
assign block_a_halt_en_active = widget_if.addr == 8;
assign block_a_halt_en_sw_wr = block_a_halt_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_a_halt_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_halt_en__crc_error_q <= 1'd0;
end
else
begin
    if (block_a_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_halt_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_a_halt_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_a_halt_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_halt_en__len_error_q <= 1'd0;
end
else
begin
    if (block_a_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_halt_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_a_halt_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_a_halt_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_a_halt_en__multi_bit_ecc_error_q <= 1'd1;
end
else
begin
    if (block_a_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_a_halt_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_a_halt_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_a_halt_en_data_mux_in = {{29{1'b0}}, block_a_halt_en__multi_bit_ecc_error_q, block_a_halt_en__len_error_q, block_a_halt_en__crc_error_q};

// Internal registers are ready immediately
assign block_a_halt_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_a_halt_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_b_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_b_int_active                      ;
logic        block_b_int_sw_wr                       ;
logic [31:0] block_b_int_data_mux_in                 ;
logic        block_b_int_rdy_mux_in                  ;
logic        block_b_int_err_mux_in                  ;
logic [0:0]  block_b_int__crc_error_q                ;
logic [0:0]  block_b_int__crc_error_sticky_latch     ;
logic [0:0]  block_b_int__len_error_q                ;
logic [0:0]  block_b_int__len_error_sticky_latch     ;
logic [0:0]  block_b_int__multi_bit_ecc_error_q      ;
logic [0:0]  block_b_int__multi_bit_ecc_error_sticky_latch;
logic [3:0]  block_b_int__active_ecc_master_q        ;
logic [3:0]  block_b_int__active_ecc_master_sticky_latch;


// Register-activation for 'block_b_int' 
assign block_b_int_active = widget_if.addr == 256;
assign block_b_int_sw_wr = block_b_int_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_b_int[0:0])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int__crc_error_q <= 1'd0;
end
else
begin
    if (block_b_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_b_int__crc_error_q[0:0] <= block_b_int__crc_error_q[0:0] & ~widget_if.w_data[0:0];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_b_int__crc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_b_int__crc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_b_int__crc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_b_int__crc_error_sticky_latch = block_b_int__crc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_b_int[1:1])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int__len_error_q <= 1'd0;
end
else
begin
    if (block_b_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_b_int__len_error_q[0:0] <= block_b_int__len_error_q[0:0] & ~widget_if.w_data[1:1];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_b_int__len_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_b_int__len_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_b_int__len_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_b_int__len_error_sticky_latch = block_b_int__len_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_b_int[2:2])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_b_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_b_int__multi_bit_ecc_error_q[0:0] <= block_b_int__multi_bit_ecc_error_q[0:0] & ~widget_if.w_data[2:2];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_b_int__multi_bit_ecc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_b_int__multi_bit_ecc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_b_int__multi_bit_ecc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_b_int__multi_bit_ecc_error_sticky_latch = block_b_int__multi_bit_ecc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : active_ecc_master (block_b_int[7:4])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'sticky']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int__active_ecc_master_q <= 4'd0;
end
else
begin
    if (block_b_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_b_int__active_ecc_master_q[3:0] <= block_b_int__active_ecc_master_q[3:0] & ~widget_if.w_data[7:4];
        end
    end
    else
    if (|block_b_int__active_ecc_master_sticky_latch && !(|block_b_int__active_ecc_master_q))
    begin
        // Sticky. Keep value until software clears it
        block_b_int__active_ecc_master_q <= block_b_int__active_ecc_master_in;
    end
end // of block_b_int__active_ecc_master's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_b_int__active_ecc_master_sticky_latch = block_b_int__active_ecc_master_in;


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign block_b_int_intr = |(block_b_int__crc_error_q & block_b_int_en__crc_error_q) || |(block_b_int__len_error_q & block_b_int_en__len_error_q) || |(block_b_int__multi_bit_ecc_error_q & block_b_int_en__multi_bit_ecc_error_q);

// Register has at least one interrupt field with halt property set
assign block_b_int_halt = |(block_b_int__crc_error_q & ~block_b_halt_en__crc_error_q) || |(block_b_int__len_error_q & ~block_b_halt_en__len_error_q) || |(block_b_int__multi_bit_ecc_error_q & ~block_b_halt_en__multi_bit_ecc_error_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_b_int_data_mux_in = {{24{1'b0}}, block_b_int__active_ecc_master_q, {1{1'b0}}, block_b_int__multi_bit_ecc_error_q, block_b_int__len_error_q, block_b_int__crc_error_q};

// Internal registers are ready immediately
assign block_b_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_b_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_b_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_b_int_en_active                ;
logic        block_b_int_en_sw_wr                 ;
logic [31:0] block_b_int_en_data_mux_in           ;
logic        block_b_int_en_rdy_mux_in            ;
logic        block_b_int_en_err_mux_in            ;
logic [0:0]  block_b_int_en__crc_error_q          ;
logic [0:0]  block_b_int_en__len_error_q          ;
logic [0:0]  block_b_int_en__multi_bit_ecc_error_q;


// Register-activation for 'block_b_int_en' 
assign block_b_int_en_active = widget_if.addr == 260;
assign block_b_int_en_sw_wr = block_b_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_b_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int_en__crc_error_q <= 1'd1;
end
else
begin
    if (block_b_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_int_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_b_int_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_b_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int_en__len_error_q <= 1'd1;
end
else
begin
    if (block_b_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_int_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_b_int_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_b_int_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_int_en__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_b_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_int_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_b_int_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_b_int_en_data_mux_in = {{29{1'b0}}, block_b_int_en__multi_bit_ecc_error_q, block_b_int_en__len_error_q, block_b_int_en__crc_error_q};

// Internal registers are ready immediately
assign block_b_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_b_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_b_halt_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_b_halt_en_active                ;
logic        block_b_halt_en_sw_wr                 ;
logic [31:0] block_b_halt_en_data_mux_in           ;
logic        block_b_halt_en_rdy_mux_in            ;
logic        block_b_halt_en_err_mux_in            ;
logic [0:0]  block_b_halt_en__crc_error_q          ;
logic [0:0]  block_b_halt_en__len_error_q          ;
logic [0:0]  block_b_halt_en__multi_bit_ecc_error_q;


// Register-activation for 'block_b_halt_en' 
assign block_b_halt_en_active = widget_if.addr == 264;
assign block_b_halt_en_sw_wr = block_b_halt_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_b_halt_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_halt_en__crc_error_q <= 1'd0;
end
else
begin
    if (block_b_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_halt_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_b_halt_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_b_halt_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_halt_en__len_error_q <= 1'd0;
end
else
begin
    if (block_b_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_halt_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_b_halt_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_b_halt_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_b_halt_en__multi_bit_ecc_error_q <= 1'd1;
end
else
begin
    if (block_b_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_b_halt_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_b_halt_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_b_halt_en_data_mux_in = {{29{1'b0}}, block_b_halt_en__multi_bit_ecc_error_q, block_b_halt_en__len_error_q, block_b_halt_en__crc_error_q};

// Internal registers are ready immediately
assign block_b_halt_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_b_halt_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_c_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_c_int_active                      ;
logic        block_c_int_sw_wr                       ;
logic [31:0] block_c_int_data_mux_in                 ;
logic        block_c_int_rdy_mux_in                  ;
logic        block_c_int_err_mux_in                  ;
logic [0:0]  block_c_int__crc_error_q                ;
logic [0:0]  block_c_int__crc_error_sticky_latch     ;
logic [0:0]  block_c_int__len_error_q                ;
logic [0:0]  block_c_int__len_error_sticky_latch     ;
logic [0:0]  block_c_int__multi_bit_ecc_error_q      ;
logic [0:0]  block_c_int__multi_bit_ecc_error_sticky_latch;
logic [3:0]  block_c_int__active_ecc_master_q        ;
logic [3:0]  block_c_int__active_ecc_master_sticky_latch;


// Register-activation for 'block_c_int' 
assign block_c_int_active = widget_if.addr == 512;
assign block_c_int_sw_wr = block_c_int_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_c_int[0:0])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int__crc_error_q <= 1'd0;
end
else
begin
    if (block_c_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_c_int__crc_error_q[0:0] <= block_c_int__crc_error_q[0:0] & ~widget_if.w_data[0:0];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_c_int__crc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_c_int__crc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_c_int__crc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_c_int__crc_error_sticky_latch = block_c_int__crc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_c_int[1:1])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int__len_error_q <= 1'd0;
end
else
begin
    if (block_c_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_c_int__len_error_q[0:0] <= block_c_int__len_error_q[0:0] & ~widget_if.w_data[1:1];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_c_int__len_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_c_int__len_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_c_int__len_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_c_int__len_error_sticky_latch = block_c_int__len_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_c_int[2:2])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_c_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_c_int__multi_bit_ecc_error_q[0:0] <= block_c_int__multi_bit_ecc_error_q[0:0] & ~widget_if.w_data[2:2];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_c_int__multi_bit_ecc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_c_int__multi_bit_ecc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_c_int__multi_bit_ecc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_c_int__multi_bit_ecc_error_sticky_latch = block_c_int__multi_bit_ecc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : active_ecc_master (block_c_int[7:4])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'sticky']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int__active_ecc_master_q <= 4'd0;
end
else
begin
    if (block_c_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_c_int__active_ecc_master_q[3:0] <= block_c_int__active_ecc_master_q[3:0] & ~widget_if.w_data[7:4];
        end
    end
    else
    if (|block_c_int__active_ecc_master_sticky_latch && !(|block_c_int__active_ecc_master_q))
    begin
        // Sticky. Keep value until software clears it
        block_c_int__active_ecc_master_q <= block_c_int__active_ecc_master_in;
    end
end // of block_c_int__active_ecc_master's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_c_int__active_ecc_master_sticky_latch = block_c_int__active_ecc_master_in;


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign block_c_int_intr = |(block_c_int__crc_error_q & block_c_int_en__crc_error_q) || |(block_c_int__len_error_q & block_c_int_en__len_error_q) || |(block_c_int__multi_bit_ecc_error_q & block_c_int_en__multi_bit_ecc_error_q);

// Register has at least one interrupt field with halt property set
assign block_c_int_halt = |(block_c_int__crc_error_q & ~block_c_halt_en__crc_error_q) || |(block_c_int__len_error_q & ~block_c_halt_en__len_error_q) || |(block_c_int__multi_bit_ecc_error_q & ~block_c_halt_en__multi_bit_ecc_error_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_c_int_data_mux_in = {{24{1'b0}}, block_c_int__active_ecc_master_q, {1{1'b0}}, block_c_int__multi_bit_ecc_error_q, block_c_int__len_error_q, block_c_int__crc_error_q};

// Internal registers are ready immediately
assign block_c_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_c_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_c_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_c_int_en_active                ;
logic        block_c_int_en_sw_wr                 ;
logic [31:0] block_c_int_en_data_mux_in           ;
logic        block_c_int_en_rdy_mux_in            ;
logic        block_c_int_en_err_mux_in            ;
logic [0:0]  block_c_int_en__crc_error_q          ;
logic [0:0]  block_c_int_en__len_error_q          ;
logic [0:0]  block_c_int_en__multi_bit_ecc_error_q;


// Register-activation for 'block_c_int_en' 
assign block_c_int_en_active = widget_if.addr == 516;
assign block_c_int_en_sw_wr = block_c_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_c_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int_en__crc_error_q <= 1'd1;
end
else
begin
    if (block_c_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_int_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_c_int_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_c_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int_en__len_error_q <= 1'd1;
end
else
begin
    if (block_c_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_int_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_c_int_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_c_int_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_int_en__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_c_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_int_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_c_int_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_c_int_en_data_mux_in = {{29{1'b0}}, block_c_int_en__multi_bit_ecc_error_q, block_c_int_en__len_error_q, block_c_int_en__crc_error_q};

// Internal registers are ready immediately
assign block_c_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_c_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_c_halt_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_c_halt_en_active                ;
logic        block_c_halt_en_sw_wr                 ;
logic [31:0] block_c_halt_en_data_mux_in           ;
logic        block_c_halt_en_rdy_mux_in            ;
logic        block_c_halt_en_err_mux_in            ;
logic [0:0]  block_c_halt_en__crc_error_q          ;
logic [0:0]  block_c_halt_en__len_error_q          ;
logic [0:0]  block_c_halt_en__multi_bit_ecc_error_q;


// Register-activation for 'block_c_halt_en' 
assign block_c_halt_en_active = widget_if.addr == 520;
assign block_c_halt_en_sw_wr = block_c_halt_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_c_halt_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_halt_en__crc_error_q <= 1'd0;
end
else
begin
    if (block_c_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_halt_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_c_halt_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_c_halt_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_halt_en__len_error_q <= 1'd0;
end
else
begin
    if (block_c_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_halt_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_c_halt_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_c_halt_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_c_halt_en__multi_bit_ecc_error_q <= 1'd1;
end
else
begin
    if (block_c_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_c_halt_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_c_halt_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_c_halt_en_data_mux_in = {{29{1'b0}}, block_c_halt_en__multi_bit_ecc_error_q, block_c_halt_en__len_error_q, block_c_halt_en__crc_error_q};

// Internal registers are ready immediately
assign block_c_halt_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_c_halt_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_d_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_d_int_active                      ;
logic        block_d_int_sw_wr                       ;
logic [31:0] block_d_int_data_mux_in                 ;
logic        block_d_int_rdy_mux_in                  ;
logic        block_d_int_err_mux_in                  ;
logic [0:0]  block_d_int__crc_error_q                ;
logic [0:0]  block_d_int__crc_error_sticky_latch     ;
logic [0:0]  block_d_int__len_error_q                ;
logic [0:0]  block_d_int__len_error_sticky_latch     ;
logic [0:0]  block_d_int__multi_bit_ecc_error_q      ;
logic [0:0]  block_d_int__multi_bit_ecc_error_sticky_latch;
logic [3:0]  block_d_int__active_ecc_master_q        ;
logic [3:0]  block_d_int__active_ecc_master_sticky_latch;


// Register-activation for 'block_d_int' 
assign block_d_int_active = widget_if.addr == 768;
assign block_d_int_sw_wr = block_d_int_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_d_int[0:0])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int__crc_error_q <= 1'd0;
end
else
begin
    if (block_d_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_d_int__crc_error_q[0:0] <= block_d_int__crc_error_q[0:0] & ~widget_if.w_data[0:0];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_d_int__crc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_d_int__crc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_d_int__crc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_d_int__crc_error_sticky_latch = block_d_int__crc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_d_int[1:1])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int__len_error_q <= 1'd0;
end
else
begin
    if (block_d_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_d_int__len_error_q[0:0] <= block_d_int__len_error_q[0:0] & ~widget_if.w_data[1:1];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_d_int__len_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_d_int__len_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_d_int__len_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_d_int__len_error_sticky_latch = block_d_int__len_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_d_int[2:2])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'intr', 'intr type', 'enable', 'haltenable']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_d_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_d_int__multi_bit_ecc_error_q[0:0] <= block_d_int__multi_bit_ecc_error_q[0:0] & ~widget_if.w_data[2:2];
        end
    end
    else
    begin
        for (int i = 0; i < 1; i++)
        begin
            if (block_d_int__multi_bit_ecc_error_sticky_latch[i])
            begin
                // Stickybit. Keep value until software clears it
                block_d_int__multi_bit_ecc_error_q[i] <= 1'b1;
            end
        end
    end
end // of block_d_int__multi_bit_ecc_error's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_d_int__multi_bit_ecc_error_sticky_latch = block_d_int__multi_bit_ecc_error_in;



//-----------------FIELD SUMMARY-----------------
// name         : active_ecc_master (block_d_int[7:4])
// access       : hw = w  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'woclr', 'desc', 'sticky']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int__active_ecc_master_q <= 4'd0;
end
else
begin
    if (block_d_int_sw_wr)
    begin
        if (widget_if.byte_en[0]) // woclr property
        begin
            block_d_int__active_ecc_master_q[3:0] <= block_d_int__active_ecc_master_q[3:0] & ~widget_if.w_data[7:4];
        end
    end
    else
    if (|block_d_int__active_ecc_master_sticky_latch && !(|block_d_int__active_ecc_master_q))
    begin
        // Sticky. Keep value until software clears it
        block_d_int__active_ecc_master_q <= block_d_int__active_ecc_master_in;
    end
end // of block_d_int__active_ecc_master's always_ff

// Define signal that causes the interrupt to be set (level-type interrupt)
assign block_d_int__active_ecc_master_sticky_latch = block_d_int__active_ecc_master_in;


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign block_d_int_intr = |(block_d_int__crc_error_q & block_d_int_en__crc_error_q) || |(block_d_int__len_error_q & block_d_int_en__len_error_q) || |(block_d_int__multi_bit_ecc_error_q & block_d_int_en__multi_bit_ecc_error_q);

// Register has at least one interrupt field with halt property set
assign block_d_int_halt = |(block_d_int__crc_error_q & ~block_d_halt_en__crc_error_q) || |(block_d_int__len_error_q & ~block_d_halt_en__len_error_q) || |(block_d_int__multi_bit_ecc_error_q & ~block_d_halt_en__multi_bit_ecc_error_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_d_int_data_mux_in = {{24{1'b0}}, block_d_int__active_ecc_master_q, {1{1'b0}}, block_d_int__multi_bit_ecc_error_q, block_d_int__len_error_q, block_d_int__crc_error_q};

// Internal registers are ready immediately
assign block_d_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_d_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_d_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_d_int_en_active                ;
logic        block_d_int_en_sw_wr                 ;
logic [31:0] block_d_int_en_data_mux_in           ;
logic        block_d_int_en_rdy_mux_in            ;
logic        block_d_int_en_err_mux_in            ;
logic [0:0]  block_d_int_en__crc_error_q          ;
logic [0:0]  block_d_int_en__len_error_q          ;
logic [0:0]  block_d_int_en__multi_bit_ecc_error_q;


// Register-activation for 'block_d_int_en' 
assign block_d_int_en_active = widget_if.addr == 772;
assign block_d_int_en_sw_wr = block_d_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_d_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int_en__crc_error_q <= 1'd1;
end
else
begin
    if (block_d_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_int_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_d_int_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_d_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int_en__len_error_q <= 1'd1;
end
else
begin
    if (block_d_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_int_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_d_int_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_d_int_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_int_en__multi_bit_ecc_error_q <= 1'd0;
end
else
begin
    if (block_d_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_int_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_d_int_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_d_int_en_data_mux_in = {{29{1'b0}}, block_d_int_en__multi_bit_ecc_error_q, block_d_int_en__len_error_q, block_d_int_en__crc_error_q};

// Internal registers are ready immediately
assign block_d_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_d_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : block_d_halt_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        block_d_halt_en_active                ;
logic        block_d_halt_en_sw_wr                 ;
logic [31:0] block_d_halt_en_data_mux_in           ;
logic        block_d_halt_en_rdy_mux_in            ;
logic        block_d_halt_en_err_mux_in            ;
logic [0:0]  block_d_halt_en__crc_error_q          ;
logic [0:0]  block_d_halt_en__len_error_q          ;
logic [0:0]  block_d_halt_en__multi_bit_ecc_error_q;


// Register-activation for 'block_d_halt_en' 
assign block_d_halt_en_active = widget_if.addr == 776;
assign block_d_halt_en_sw_wr = block_d_halt_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : crc_error (block_d_halt_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_halt_en__crc_error_q <= 1'd0;
end
else
begin
    if (block_d_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_halt_en__crc_error_q[0:0] <= widget_if.w_data[0:0];
    end
end // of block_d_halt_en__crc_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : len_error (block_d_halt_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_halt_en__len_error_q <= 1'd0;
end
else
begin
    if (block_d_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_halt_en__len_error_q[0:0] <= widget_if.w_data[1:1];
    end
end // of block_d_halt_en__len_error's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : multi_bit_ecc_error (block_d_halt_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    block_d_halt_en__multi_bit_ecc_error_q <= 1'd1;
end
else
begin
    if (block_d_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            block_d_halt_en__multi_bit_ecc_error_q[0:0] <= widget_if.w_data[2:2];
    end
end // of block_d_halt_en__multi_bit_ecc_error's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign block_d_halt_en_data_mux_in = {{29{1'b0}}, block_d_halt_en__multi_bit_ecc_error_q, block_d_halt_en__len_error_q, block_d_halt_en__crc_error_q};

// Internal registers are ready immediately
assign block_d_halt_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign block_d_halt_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : master_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        master_int_active         ;
logic [31:0] master_int_data_mux_in    ;
logic        master_int_rdy_mux_in     ;
logic        master_int_err_mux_in     ;
logic [0:0]  master_int__module_a_int_q;
logic [0:0]  master_int__module_b_int_q;
logic [0:0]  master_int__module_c_int_q;
logic [0:0]  master_int__module_d_int_q;


// Register-activation for 'master_int' 
assign master_int_active = widget_if.addr == 4096;

//-----------------FIELD SUMMARY-----------------
// name         : module_a_int (master_int[0:0])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'enable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int__module_a_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_int__module_a_int_q <= block_a_int_intr;
    end
end // of master_int__module_a_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_b_int (master_int[1:1])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'enable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int__module_b_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_int__module_b_int_q <= block_b_int_intr;
    end
end // of master_int__module_b_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_c_int (master_int[2:2])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'enable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int__module_c_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_int__module_c_int_q <= block_c_int_intr;
    end
end // of master_int__module_c_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_d_int (master_int[3:3])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'enable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int__module_d_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_int__module_d_int_q <= block_d_int_intr;
    end
end // of master_int__module_d_int's always_ff


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign master_int_intr = |(master_int__module_a_int_q & master_int_en__module_a_int_en_q) || |(master_int__module_b_int_q & master_int_en__module_b_int_en_q) || |(master_int__module_c_int_q & master_int_en__module_c_int_en_q) || |(master_int__module_d_int_q & master_int_en__module_d_int_en_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign master_int_data_mux_in = {{28{1'b0}}, master_int__module_d_int_q, master_int__module_c_int_q, master_int__module_b_int_q, master_int__module_a_int_q};

// Internal registers are ready immediately
assign master_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign master_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (1'b0)));

/*******************************************************************
/*******************************************************************
/* REGISTER              : master_halt
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        master_halt_active         ;
logic [31:0] master_halt_data_mux_in    ;
logic        master_halt_rdy_mux_in     ;
logic        master_halt_err_mux_in     ;
logic [0:0]  master_halt__module_a_int_q;
logic [0:0]  master_halt__module_b_int_q;
logic [0:0]  master_halt__module_c_int_q;
logic [0:0]  master_halt__module_d_int_q;


// Register-activation for 'master_halt' 
assign master_halt_active = widget_if.addr == 4100;

//-----------------FIELD SUMMARY-----------------
// name         : module_a_int (master_halt[0:0])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'haltenable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt__module_a_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_halt__module_a_int_q <= block_a_int_halt;
    end
end // of master_halt__module_a_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_b_int (master_halt[1:1])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'haltenable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt__module_b_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_halt__module_b_int_q <= block_b_int_halt;
    end
end // of master_halt__module_b_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_c_int (master_halt[2:2])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'haltenable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt__module_c_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_halt__module_c_int_q <= block_c_int_halt;
    end
end // of master_halt__module_c_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_d_int (master_halt[3:3])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['intr', 'stickybit', 'sw', 'desc', 'haltenable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt__module_d_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        master_halt__module_d_int_q <= block_d_int_halt;
    end
end // of master_halt__module_d_int's always_ff


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign master_halt_intr = |(master_halt__module_a_int_q) || |(master_halt__module_b_int_q) || |(master_halt__module_c_int_q) || |(master_halt__module_d_int_q);

// Register has at least one interrupt field with halt property set
assign master_halt_halt = |(master_halt__module_a_int_q & ~master_halt_en__module_a_halt_en_q) || |(master_halt__module_b_int_q & ~master_halt_en__module_b_halt_en_q) || |(master_halt__module_c_int_q & ~master_halt_en__module_c_halt_en_q) || |(master_halt__module_d_int_q & ~master_halt_en__module_d_halt_en_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign master_halt_data_mux_in = {{28{1'b0}}, master_halt__module_d_int_q, master_halt__module_c_int_q, master_halt__module_b_int_q, master_halt__module_a_int_q};

// Internal registers are ready immediately
assign master_halt_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign master_halt_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (1'b0)));

/*******************************************************************
/*******************************************************************
/* REGISTER              : master_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        master_int_en_active            ;
logic        master_int_en_sw_wr             ;
logic [31:0] master_int_en_data_mux_in       ;
logic        master_int_en_rdy_mux_in        ;
logic        master_int_en_err_mux_in        ;
logic [0:0]  master_int_en__module_a_int_en_q;
logic [0:0]  master_int_en__module_b_int_en_q;
logic [0:0]  master_int_en__module_c_int_en_q;
logic [0:0]  master_int_en__module_d_int_en_q;


// Register-activation for 'master_int_en' 
assign master_int_en_active = widget_if.addr == 4104;
assign master_int_en_sw_wr = master_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : module_a_int_en (master_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int_en__module_a_int_en_q <= 1'd0;
end
else
begin
    if (master_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_int_en__module_a_int_en_q[0:0] <= widget_if.w_data[0:0];
    end
end // of master_int_en__module_a_int_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_b_int_en (master_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int_en__module_b_int_en_q <= 1'd0;
end
else
begin
    if (master_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_int_en__module_b_int_en_q[0:0] <= widget_if.w_data[1:1];
    end
end // of master_int_en__module_b_int_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_c_int_en (master_int_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int_en__module_c_int_en_q <= 1'd0;
end
else
begin
    if (master_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_int_en__module_c_int_en_q[0:0] <= widget_if.w_data[2:2];
    end
end // of master_int_en__module_c_int_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_d_int_en (master_int_en[3:3])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_int_en__module_d_int_en_q <= 1'd0;
end
else
begin
    if (master_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_int_en__module_d_int_en_q[0:0] <= widget_if.w_data[3:3];
    end
end // of master_int_en__module_d_int_en's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign master_int_en_data_mux_in = {{28{1'b0}}, master_int_en__module_d_int_en_q, master_int_en__module_c_int_en_q, master_int_en__module_b_int_en_q, master_int_en__module_a_int_en_q};

// Internal registers are ready immediately
assign master_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign master_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : master_halt_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        master_halt_en_active             ;
logic        master_halt_en_sw_wr              ;
logic [31:0] master_halt_en_data_mux_in        ;
logic        master_halt_en_rdy_mux_in         ;
logic        master_halt_en_err_mux_in         ;
logic [0:0]  master_halt_en__module_a_halt_en_q;
logic [0:0]  master_halt_en__module_b_halt_en_q;
logic [0:0]  master_halt_en__module_c_halt_en_q;
logic [0:0]  master_halt_en__module_d_halt_en_q;


// Register-activation for 'master_halt_en' 
assign master_halt_en_active = widget_if.addr == 4108;
assign master_halt_en_sw_wr = master_halt_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : module_a_halt_en (master_halt_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt_en__module_a_halt_en_q <= 1'd0;
end
else
begin
    if (master_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_halt_en__module_a_halt_en_q[0:0] <= widget_if.w_data[0:0];
    end
end // of master_halt_en__module_a_halt_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_b_halt_en (master_halt_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt_en__module_b_halt_en_q <= 1'd0;
end
else
begin
    if (master_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_halt_en__module_b_halt_en_q[0:0] <= widget_if.w_data[1:1];
    end
end // of master_halt_en__module_b_halt_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_c_halt_en (master_halt_en[2:2])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt_en__module_c_halt_en_q <= 1'd0;
end
else
begin
    if (master_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_halt_en__module_c_halt_en_q[0:0] <= widget_if.w_data[2:2];
    end
end // of master_halt_en__module_c_halt_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : module_d_halt_en (master_halt_en[3:3])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    master_halt_en__module_d_halt_en_q <= 1'd0;
end
else
begin
    if (master_halt_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            master_halt_en__module_d_halt_en_q[0:0] <= widget_if.w_data[3:3];
    end
end // of master_halt_en__module_d_halt_en's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign master_halt_en_data_mux_in = {{28{1'b0}}, master_halt_en__module_d_halt_en_q, master_halt_en__module_c_halt_en_q, master_halt_en__module_b_halt_en_q, master_halt_en__module_a_halt_en_q};

// Internal registers are ready immediately
assign master_halt_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign master_halt_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

/*******************************************************************
/*******************************************************************
/* REGISTER              : global_int
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        global_int_active        ;
logic [31:0] global_int_data_mux_in   ;
logic        global_int_rdy_mux_in    ;
logic        global_int_err_mux_in    ;
logic [0:0]  global_int__global_int_q ;
logic [0:0]  global_int__global_halt_q;


// Register-activation for 'global_int' 
assign global_int_active = widget_if.addr == 4112;

//-----------------FIELD SUMMARY-----------------
// name         : global_int (global_int[0:0])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'intr', 'stickybit', 'desc', 'enable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    global_int__global_int_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        global_int__global_int_q <= master_int_intr;
    end
end // of global_int__global_int's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : global_halt (global_int[1:1])
// access       : hw = w  
//                sw = r (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'intr', 'stickybit', 'desc', 'haltenable', 'next']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    global_int__global_halt_q <= 1'd0;
end
else
begin
    begin
        // Non-sticky interrupt. Only keep value high if source keeps up
        global_int__global_halt_q <= master_halt_halt;
    end
end // of global_int__global_halt's always_ff


/************************************** 
 * Register contains interrupts    *
 **************************************/
// Register has at least one interrupt field
assign global_int_intr = |(global_int__global_int_q & global_int_en__global_int_en_q) || |(global_int__global_halt_q);

// Register has at least one interrupt field with halt property set
assign global_int_halt = |(global_int__global_int_q) || |(global_int__global_halt_q & ~global_int_en__global_halt_en_q);


/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign global_int_data_mux_in = {{30{1'b0}}, global_int__global_halt_q, global_int__global_int_q};

// Internal registers are ready immediately
assign global_int_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign global_int_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (1'b0)));

/*******************************************************************
/*******************************************************************
/* REGISTER              : global_int_en
/* DIMENSION             : 0
/* DEPTHS (per dimension): []
/*******************************************************************
/*******************************************************************/

logic        global_int_en_active           ;
logic        global_int_en_sw_wr            ;
logic [31:0] global_int_en_data_mux_in      ;
logic        global_int_en_rdy_mux_in       ;
logic        global_int_en_err_mux_in       ;
logic [0:0]  global_int_en__global_int_en_q ;
logic [0:0]  global_int_en__global_halt_en_q;


// Register-activation for 'global_int_en' 
assign global_int_en_active = widget_if.addr == 4116;
assign global_int_en_sw_wr = global_int_en_active && widget_if.w_vld;

//-----------------FIELD SUMMARY-----------------
// name         : global_int_en (global_int_en[0:0])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    global_int_en__global_int_en_q <= 1'd0;
end
else
begin
    if (global_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            global_int_en__global_int_en_q[0:0] <= widget_if.w_data[0:0];
    end
end // of global_int_en__global_int_en's always_ff



//-----------------FIELD SUMMARY-----------------
// name         : global_halt_en (global_int_en[1:1])
// access       : hw = na  
//                sw = rw (precedence)
// reset        : active_low / asynchronous
// flags        : ['sw', 'desc']
// external     : False
// storage type : StorageType.FLOPS
//-----------------------------------------------

always_ff @(posedge clk or negedge field_reset_n)
if (!field_reset_n)
begin
    global_int_en__global_halt_en_q <= 1'd0;
end
else
begin
    if (global_int_en_sw_wr)
    begin
        if (widget_if.byte_en[0])
            global_int_en__global_halt_en_q[0:0] <= widget_if.w_data[1:1];
    end
end // of global_int_en__global_halt_en's always_ff




/************************************** 
 * Assign all fields to signal to Mux *
 **************************************/
// Assign all fields. Fields that are not readable are tied to 0.
assign global_int_en_data_mux_in = {{30{1'b0}}, global_int_en__global_halt_en_q, global_int_en__global_int_en_q};

// Internal registers are ready immediately
assign global_int_en_rdy_mux_in = 1'b1;

// Return an error if *no* read and *no* write was succesful. If some bits
// cannot be read/written but others are succesful, don't return and error
// Hence, as long as one action can be succesful, no error will be returned.
assign global_int_en_err_mux_in = !((widget_if.r_vld && (widget_if.byte_en[0])) || (widget_if.w_vld && (widget_if.byte_en[0])));

// Read multiplexer
always_comb
begin
    unique case (1'b1)
        block_a_int_active:
        begin
            widget_if.r_data = block_a_int_data_mux_in;
            widget_if.err    = block_a_int_err_mux_in;
            widget_if.rdy    = block_a_int_rdy_mux_in;
        end
        block_a_int_en_active:
        begin
            widget_if.r_data = block_a_int_en_data_mux_in;
            widget_if.err    = block_a_int_en_err_mux_in;
            widget_if.rdy    = block_a_int_en_rdy_mux_in;
        end
        block_a_halt_en_active:
        begin
            widget_if.r_data = block_a_halt_en_data_mux_in;
            widget_if.err    = block_a_halt_en_err_mux_in;
            widget_if.rdy    = block_a_halt_en_rdy_mux_in;
        end
        block_b_int_active:
        begin
            widget_if.r_data = block_b_int_data_mux_in;
            widget_if.err    = block_b_int_err_mux_in;
            widget_if.rdy    = block_b_int_rdy_mux_in;
        end
        block_b_int_en_active:
        begin
            widget_if.r_data = block_b_int_en_data_mux_in;
            widget_if.err    = block_b_int_en_err_mux_in;
            widget_if.rdy    = block_b_int_en_rdy_mux_in;
        end
        block_b_halt_en_active:
        begin
            widget_if.r_data = block_b_halt_en_data_mux_in;
            widget_if.err    = block_b_halt_en_err_mux_in;
            widget_if.rdy    = block_b_halt_en_rdy_mux_in;
        end
        block_c_int_active:
        begin
            widget_if.r_data = block_c_int_data_mux_in;
            widget_if.err    = block_c_int_err_mux_in;
            widget_if.rdy    = block_c_int_rdy_mux_in;
        end
        block_c_int_en_active:
        begin
            widget_if.r_data = block_c_int_en_data_mux_in;
            widget_if.err    = block_c_int_en_err_mux_in;
            widget_if.rdy    = block_c_int_en_rdy_mux_in;
        end
        block_c_halt_en_active:
        begin
            widget_if.r_data = block_c_halt_en_data_mux_in;
            widget_if.err    = block_c_halt_en_err_mux_in;
            widget_if.rdy    = block_c_halt_en_rdy_mux_in;
        end
        block_d_int_active:
        begin
            widget_if.r_data = block_d_int_data_mux_in;
            widget_if.err    = block_d_int_err_mux_in;
            widget_if.rdy    = block_d_int_rdy_mux_in;
        end
        block_d_int_en_active:
        begin
            widget_if.r_data = block_d_int_en_data_mux_in;
            widget_if.err    = block_d_int_en_err_mux_in;
            widget_if.rdy    = block_d_int_en_rdy_mux_in;
        end
        block_d_halt_en_active:
        begin
            widget_if.r_data = block_d_halt_en_data_mux_in;
            widget_if.err    = block_d_halt_en_err_mux_in;
            widget_if.rdy    = block_d_halt_en_rdy_mux_in;
        end
        master_int_active:
        begin
            widget_if.r_data = master_int_data_mux_in;
            widget_if.err    = master_int_err_mux_in;
            widget_if.rdy    = master_int_rdy_mux_in;
        end
        master_halt_active:
        begin
            widget_if.r_data = master_halt_data_mux_in;
            widget_if.err    = master_halt_err_mux_in;
            widget_if.rdy    = master_halt_rdy_mux_in;
        end
        master_int_en_active:
        begin
            widget_if.r_data = master_int_en_data_mux_in;
            widget_if.err    = master_int_en_err_mux_in;
            widget_if.rdy    = master_int_en_rdy_mux_in;
        end
        master_halt_en_active:
        begin
            widget_if.r_data = master_halt_en_data_mux_in;
            widget_if.err    = master_halt_en_err_mux_in;
            widget_if.rdy    = master_halt_en_rdy_mux_in;
        end
        global_int_active:
        begin
            widget_if.r_data = global_int_data_mux_in;
            widget_if.err    = global_int_err_mux_in;
            widget_if.rdy    = global_int_rdy_mux_in;
        end
        global_int_en_active:
        begin
            widget_if.r_data = global_int_en_data_mux_in;
            widget_if.err    = global_int_en_err_mux_in;
            widget_if.rdy    = global_int_en_rdy_mux_in;
        end
        default:
        begin
            // If the address is not found, return an error
            widget_if.r_data = 0;
            widget_if.err    = 1;
            widget_if.rdy    = widget_if.r_vld || widget_if.w_vld;
        end
    endcase
end
endmodule
